SCHMITT CKT - ECL COMPATIBLE SCHMITT TRIGGER
.MODEL QSTD NPN
+ is=1E-14 BF=50 BR=0.1 RB=50 RC=10 TF=0.12N
+   TR=5NS CJE=0.4P VJE=0.8 MJE=0.4 CJC=0.5P VJC=0.8 MJC=0.333
+   VAF=50

RIN 1 2 50
RC1 8 3 50
R1 3 5 185
R2 5 0 760
RC2 8 6 100
RE 4 0 260
RTH1 7 0 125
RTH2 7 0 85
CLOAD 7 0 5P
Q1 3 2 4 0 QSTD
Q2 6 5 4 0 QSTD
Q3 8 6 7 0 QSTD
Q4 8 6 7 0 QSTD


VCC 8 0 5.0
VIN 1 0 pwl( 0.0ns 3.4 200ns 3.8 400ns 3.4 600ns 3.8 800ns 3.4 )

*.print tran v(1) v(6) v(7)
*.tran 1ns 500ns
.option acct limpts=1000
.op 
.end 
