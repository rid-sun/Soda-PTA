THMT9 NINE SOLUTION CIRCUIT 2001.01.23 Y.INOUE
*.OPTIONS GMIN=1N
VCC 1 0 DC 1.0
*VCC 111 0 DC 1.0
*R 111 1 10K
R1 1 121 10K
Q1 3 2 1 QP
Q2 2 3 0 QN
Q53 121 5 0 QP 20 
Q35 122 3 0 QP 40
R2 1 122 10K 
Q4 5 4 1 QP
Q5 4 5 0 QN 
*Q7 2 2 1 QP
*Q8 4 4 1 QP 10
.MODEL QN NPN (IS=1F BF=100 BR=1 RC=1K RB=100)
.MODEL QP PNP (IS=1F BF=100 BR=1 RC=1K RB=100)
*.MODEL QN NPN (IS=1F BF=100 BR=1 )
*.MODEL QP PNP (IS=1F BF=100 BR=1 )
*.END

.OPTIONS DELMAX=1000ns
.op
*.gmin
.end