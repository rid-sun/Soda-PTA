TRCKT --- Four Transistor Circuit 
*
*TEST CIRCUIT (TRCKT)
*
*.OP
*
VCC VPLUS 0  DC 12
*
RC1 VPLUS T1C 4K
RC2 VPLUS T2C 4K
RT1T2 T1C T2B 30K
RT2B T2B 0 10.1K
RT12E T12E 0 500
RT2CF T2C VINMINUS 30K 
RC3 VPLUS T3C 4K
RC4 VPLUS T4C 4K
RT3T4 T3C T4B 30K
RT4B T4B 0 10.1K
RT34E T34E 0 500
RT4CF T4C V2 30K 
RT13B T13B 0 5K
V2 V2 VINMINUS DC 2
* VIN, 25:UNIEQUE SOLUTION, 10:NINE SOLUTION
VIN VINMINUS T13B DC 10
QT1 T1C T13B T12E QNPN OFF
QT2 T2C T2B T12E QNPN
QT3 T3C T13B T34E QNPN OFF
QT4 T4C T4B T34E QNPN 
.MODEL QNPN NPN (IS=1E-9 BF=49 BR=1)
*.OPTIONS ACCT LIST NOMOD 
*.END 

.OPTIONS DELMAX=1000ns
.op
*.gmin
.end
