THMT5 FIVE, SEVEN, NINE SOLUTION CIRCUIT 2001.01.23 Y.INOUE
*ITER=336
*.OP
VCC 1 0 DC 0.44
*VCC 1 0 DC 1.0
Q1 3 2 1 QP
Q2 2 3 0 QN
Q3 4 3 0 QN 10
Q4 5 4 1 QP
Q5 4 5 0 QN
Q6 6 5 0 QN 10
Q7 7 6 1 QP
Q8 6 7 0 QN
Q31 6 3 0 QN 
.MODEL QN NPN (IS=1F BF=100 BR=1 RC=1K RB=100)
.MODEL QP PNP (IS=1F BF=100 BR=1 RC=1K RB=100)
*.OPTIONS ACCT LIST NOMOD GMIN=1N
*.OPTIONS ACCT LIST NOMOD 
*.END

.OPTIONS DELMAX=1000ns
.op
*.gmin
.end
