TADEGLOW CKT
VCC 1 0 DC 12.0
RT1C 1 2 4.0K
RT1E 3 0 0.1K
RT2B 2 5 8.0K
RT1B 6 4 8.0K
RT2C 1 6 4.0K
RT2E 7 0 0.1K
D 8 6 DIODE
RT3CD 9 8 30.0K
RT3C 1 9 1.0K
RT3E 10 0 0.1K
RT3B 11 12 10.0K
RT4C 1 12 4.0K
RT4B1 1 13 10.0K
RT4B2 13 0 1.0K
QT1 2 4 3 QNPN
QT2 6 5 7 QNPN
QT3 9 11 10 QNPN
QT4 12 13 0 QNPN
.MODEL DIODE D (IS=1.0E-14)
.MODEL QNPN NPN (IS=1.0E-14 BF=100 VAF=50)
*.END


.OPTIONS DELMAX=1000ns
.op
*.gmin
.end 