TRISTABLE CIRCUIT SHOU&GREEN 2001.5.28
* Five Solutions
*.OP
*.OPTIONS NOMOD
*.NODESET V(4)=3.3 V(5)=3.3
VDD 1 0 DC 3.3
M1 4 2 1 1 PCH W=1.3U L=0.5U 
M2 5 3 1 1 PCH W=1.3U L=0.5U
M3 4 4 3 3 NCH W=2.8U L=0.4U
M4 5 5 2 3 NCH W=2.8U L=0.4U
M5 3 5 0 0 NCH W=1.9U L=0.4U
M6 2 4 0 0 NCH W=1.9U L=0.4U
.MODEL PCH PMOS (LEVEL=8
.MODEL NCH NMOS (LEVEL=8
*.END

.OPTIONS DELMAX=1000ns
.op
*.gmin
.end 