voter.sp SPICE FILE
.model nenh nmos  level = 2    vto = 0.6    pb = 0.7   cgso = 1.5e-10   cgdo = 1.5e-10    rsh = 28   cj = 0.000175    mj = 0.65   cjsw = 4e-10   mjsw = 0.3    tox = 3.5e-08   nsub = 7e+15    xj = 2e-07   ld = 2.5e-07   uo = 700    ucrit = 70000   uexp = 0.13    vmax = 50000   neff = 3    delta = 1.5
.model penh pmos  level = 2    vto = -0.6    pb = 0.7   cgso = 1.3e-10   cgdo = 1.3e-10    rsh = 92   cj = 0.000225    mj = 0.5   cjsw = 3e-10   mjsw = 0.3    tox = 3.5e-08   nsub = 5e+15    xj = 1e-07   ld = 2.5e-07   uo = 270    ucrit = 90000   uexp = 0.35    vmax = 30000   neff = 1.5    delta = 1
m1 3 5 4 3 penh l=2e-06 w=9.7e-05 

m2 4 5 3 3 penh l=2e-06 w=9.5e-05 

m3 3 5 4 3 penh l=2e-06 w=9.5e-05 

m4 4 5 3 3 penh l=2e-06 w=9.6e-05 

m5 3 5 4 3 penh l=2e-06 w=9.6e-05 

m6 4 5 3 3 penh l=2e-06 w=9.5e-05 

m7 3 5 4 3 penh l=2e-06 w=9.5e-05 

m8 4 5 3 3 penh l=2e-06 w=9.6e-05 

m9 3 6 5 3 penh l=2e-06 w=5.3e-05 

m10 5 6 3 3 penh l=2e-06 w=5.3e-05 

m11 3 7 6 3 penh l=2e-06 w=4.9e-05 

m12 7 8 3 3 penh l=2e-06 w=2.3e-05 

m13 3 6 5 3 penh l=2e-06 w=4.8e-05 

m14 5 6 3 3 penh l=2e-06 w=4.8e-05 

m15 3 8 9 3 penh l=2e-06 w=2.2e-05 

m16 10 11 3 3 penh l=2e-06 w=5e-05 

m17 3 9 11 3 penh l=2e-06 w=4.7e-05 

m18 10 11 3 3 penh l=2e-06 w=4.8e-05 

m19 3 11 10 3 penh l=2e-06 w=4.8e-05 

m20 0 10 4 0 nenh l=2e-06 w=4.6e-05 

m21 4 10 0 0 nenh l=2e-06 w=4.8e-05 

m22 0 10 4 0 nenh l=2e-06 w=4.6e-05 

m23 4 10 0 0 nenh l=2e-06 w=4.8e-05 

m24 0 10 4 0 nenh l=2e-06 w=4.8e-05 

m25 4 10 0 0 nenh l=2e-06 w=4.8e-05 

m26 0 10 4 0 nenh l=2e-06 w=4.8e-05 

m27 4 10 0 0 nenh l=2e-06 w=4.6e-05 

m28 0 11 10 0 nenh l=2e-06 w=6e-05 

m29 10 11 0 0 nenh l=2e-06 w=6e-05 

m30 11 9 0 0 nenh l=2e-06 w=5e-05 

m31 0 6 5 0 nenh l=2e-06 w=3.5e-05 

m32 5 6 0 0 nenh l=2e-06 w=3.4e-05 

m33 0 8 9 0 nenh l=2e-06 w=2.4e-05 

m34 0 6 5 0 nenh l=2e-06 w=2.5e-05 

m35 5 6 0 0 nenh l=2e-06 w=2.5e-05 

m36 0 7 6 0 nenh l=2e-06 w=1.6e-05 

m37 7 8 0 0 nenh l=2e-06 w=2.3e-05 

m38 3 13 12 3 penh l=2e-06 w=9.7e-05 

m39 12 13 3 3 penh l=2e-06 w=9.5e-05 

m40 3 13 12 3 penh l=2e-06 w=9.5e-05 

m41 12 13 3 3 penh l=2e-06 w=9.6e-05 

m42 3 13 12 3 penh l=2e-06 w=9.6e-05 

m43 12 13 3 3 penh l=2e-06 w=9.5e-05 

m44 3 13 12 3 penh l=2e-06 w=9.5e-05 

m45 12 13 3 3 penh l=2e-06 w=9.6e-05 

m46 3 14 13 3 penh l=2e-06 w=5.3e-05 

m47 13 14 3 3 penh l=2e-06 w=5.3e-05 

m48 3 15 14 3 penh l=2e-06 w=4.9e-05 

m49 15 16 3 3 penh l=2e-06 w=2.3e-05 

m50 3 14 13 3 penh l=2e-06 w=4.8e-05 

m51 13 14 3 3 penh l=2e-06 w=4.8e-05 

m52 3 16 17 3 penh l=2e-06 w=2.2e-05 

m53 18 19 3 3 penh l=2e-06 w=5e-05 

m54 3 17 19 3 penh l=2e-06 w=4.7e-05 

m55 18 19 3 3 penh l=2e-06 w=4.8e-05 

m56 3 19 18 3 penh l=2e-06 w=4.8e-05 

m57 0 18 12 0 nenh l=2e-06 w=4.6e-05 

m58 12 18 0 0 nenh l=2e-06 w=4.8e-05 

m59 0 18 12 0 nenh l=2e-06 w=4.6e-05 

m60 12 18 0 0 nenh l=2e-06 w=4.8e-05 

m61 0 18 12 0 nenh l=2e-06 w=4.8e-05 

m62 12 18 0 0 nenh l=2e-06 w=4.8e-05 

m63 0 18 12 0 nenh l=2e-06 w=4.8e-05 

m64 12 18 0 0 nenh l=2e-06 w=4.6e-05 

m65 0 19 18 0 nenh l=2e-06 w=6e-05 

m66 18 19 0 0 nenh l=2e-06 w=6e-05 

m67 19 17 0 0 nenh l=2e-06 w=5e-05 

m68 0 14 13 0 nenh l=2e-06 w=3.5e-05 

m69 13 14 0 0 nenh l=2e-06 w=3.4e-05 

m70 0 16 17 0 nenh l=2e-06 w=2.4e-05 

m71 0 14 13 0 nenh l=2e-06 w=2.5e-05 

m72 13 14 0 0 nenh l=2e-06 w=2.5e-05 

m73 0 15 14 0 nenh l=2e-06 w=1.6e-05 

m74 15 16 0 0 nenh l=2e-06 w=2.3e-05 

m75 3 21 20 3 penh l=2e-06 w=9.7e-05 

m76 20 21 3 3 penh l=2e-06 w=9.5e-05 

m77 3 21 20 3 penh l=2e-06 w=9.5e-05 

m78 20 21 3 3 penh l=2e-06 w=9.6e-05 

m79 3 21 20 3 penh l=2e-06 w=9.6e-05 

m80 20 21 3 3 penh l=2e-06 w=9.5e-05 

m81 3 21 20 3 penh l=2e-06 w=9.5e-05 

m82 20 21 3 3 penh l=2e-06 w=9.6e-05 

m83 3 22 21 3 penh l=2e-06 w=5.3e-05 

m84 21 22 3 3 penh l=2e-06 w=5.3e-05 

m85 3 23 22 3 penh l=2e-06 w=4.9e-05 

m86 23 24 3 3 penh l=2e-06 w=2.3e-05 

m87 3 22 21 3 penh l=2e-06 w=4.8e-05 

m88 21 22 3 3 penh l=2e-06 w=4.8e-05 

m89 3 24 25 3 penh l=2e-06 w=2.2e-05 

m90 26 27 3 3 penh l=2e-06 w=5e-05 

m91 3 25 27 3 penh l=2e-06 w=4.7e-05 

m92 26 27 3 3 penh l=2e-06 w=4.8e-05 

m93 3 27 26 3 penh l=2e-06 w=4.8e-05 

m94 0 26 20 0 nenh l=2e-06 w=4.6e-05 

m95 20 26 0 0 nenh l=2e-06 w=4.8e-05 

m96 0 26 20 0 nenh l=2e-06 w=4.6e-05 

m97 20 26 0 0 nenh l=2e-06 w=4.8e-05 

m98 0 26 20 0 nenh l=2e-06 w=4.8e-05 

m99 20 26 0 0 nenh l=2e-06 w=4.8e-05 

m100 0 26 20 0 nenh l=2e-06 w=4.8e-05 

m101 20 26 0 0 nenh l=2e-06 w=4.6e-05 

m102 0 27 26 0 nenh l=2e-06 w=6e-05 

m103 26 27 0 0 nenh l=2e-06 w=6e-05 

m104 27 25 0 0 nenh l=2e-06 w=5e-05 

m105 0 22 21 0 nenh l=2e-06 w=3.5e-05 

m106 21 22 0 0 nenh l=2e-06 w=3.4e-05 

m107 0 24 25 0 nenh l=2e-06 w=2.4e-05 

m108 0 22 21 0 nenh l=2e-06 w=2.5e-05 

m109 21 22 0 0 nenh l=2e-06 w=2.5e-05 

m110 0 23 22 0 nenh l=2e-06 w=1.6e-05 

m111 23 24 0 0 nenh l=2e-06 w=2.3e-05 

m112 28 29 3 3 penh l=2e-06 w=6.2e-05 

m113 3 30 29 3 penh l=2e-06 w=6.2e-05 

m114 30 31 3 3 penh l=2e-06 w=2.9e-05 

m115 3 32 31 3 penh l=4e-06 w=2.9e-05 

m116 30 31 0 0 nenh l=2e-06 w=2.1e-05 

m117 0 32 31 0 nenh l=4e-06 w=2.1e-05 

m118 28 29 0 0 nenh l=2e-06 w=4.8e-05 

m119 0 30 29 0 nenh l=2e-06 w=4.8e-05 

m120 32 0 0 0 nenh l=4e-06 w=2.5e-05 

m121 33 34 3 3 penh l=2e-06 w=6.2e-05 

m122 3 35 34 3 penh l=2e-06 w=6.2e-05 

m123 35 36 3 3 penh l=2e-06 w=2.9e-05 

m124 3 37 36 3 penh l=4e-06 w=2.9e-05 

m125 35 36 0 0 nenh l=2e-06 w=2.1e-05 

m126 0 37 36 0 nenh l=4e-06 w=2.1e-05 

m127 33 34 0 0 nenh l=2e-06 w=4.8e-05 

m128 0 35 34 0 nenh l=2e-06 w=4.8e-05 

m129 37 0 0 0 nenh l=4e-06 w=2.5e-05 

m130 38 39 3 3 penh l=2e-06 w=6.2e-05 

m131 3 40 39 3 penh l=2e-06 w=6.2e-05 

m132 40 41 3 3 penh l=2e-06 w=2.9e-05 

m133 3 42 41 3 penh l=4e-06 w=2.9e-05 

m134 40 41 0 0 nenh l=2e-06 w=2.1e-05 

m135 0 42 41 0 nenh l=4e-06 w=2.1e-05 

m136 38 39 0 0 nenh l=2e-06 w=4.8e-05 

m137 0 40 39 0 nenh l=2e-06 w=4.8e-05 

m138 42 0 0 0 nenh l=4e-06 w=2.5e-05 

m139 43 44 3 3 penh l=2e-06 w=6.2e-05 

m140 3 45 44 3 penh l=2e-06 w=6.2e-05 

m141 45 46 3 3 penh l=2e-06 w=2.9e-05 

m142 3 47 46 3 penh l=4e-06 w=2.9e-05 

m143 45 46 0 0 nenh l=2e-06 w=2.1e-05 

m144 0 47 46 0 nenh l=4e-06 w=2.1e-05 

m145 43 44 0 0 nenh l=2e-06 w=4.8e-05 

m146 0 45 44 0 nenh l=2e-06 w=4.8e-05 

m147 47 0 0 0 nenh l=4e-06 w=2.5e-05 

m148 48 49 3 3 penh l=2e-06 w=6.2e-05 

m149 3 50 49 3 penh l=2e-06 w=6.2e-05 

m150 50 51 3 3 penh l=2e-06 w=2.9e-05 

m151 3 52 51 3 penh l=4e-06 w=2.9e-05 

m152 50 51 0 0 nenh l=2e-06 w=2.1e-05 

m153 0 52 51 0 nenh l=4e-06 w=2.1e-05 

m154 48 49 0 0 nenh l=2e-06 w=4.8e-05 

m155 0 50 49 0 nenh l=2e-06 w=4.8e-05 

m156 52 0 0 0 nenh l=4e-06 w=2.5e-05 

m157 53 54 3 3 penh l=2e-06 w=6.2e-05 

m158 3 55 54 3 penh l=2e-06 w=6.2e-05 

m159 55 56 3 3 penh l=2e-06 w=2.9e-05 

m160 3 57 56 3 penh l=4e-06 w=2.9e-05 

m161 55 56 0 0 nenh l=2e-06 w=2.1e-05 

m162 0 57 56 0 nenh l=4e-06 w=2.1e-05 

m163 53 54 0 0 nenh l=2e-06 w=4.8e-05 

m164 0 55 54 0 nenh l=2e-06 w=4.8e-05 

m165 57 0 0 0 nenh l=4e-06 w=2.5e-05 

m166 3 59 58 3 penh l=2e-06 w=9.7e-05 

m167 58 59 3 3 penh l=2e-06 w=9.5e-05 

m168 3 59 58 3 penh l=2e-06 w=9.5e-05 

m169 58 59 3 3 penh l=2e-06 w=9.6e-05 

m170 3 59 58 3 penh l=2e-06 w=9.6e-05 

m171 58 59 3 3 penh l=2e-06 w=9.5e-05 

m172 3 59 58 3 penh l=2e-06 w=9.5e-05 

m173 58 59 3 3 penh l=2e-06 w=9.6e-05 

m174 3 60 59 3 penh l=2e-06 w=5.3e-05 

m175 59 60 3 3 penh l=2e-06 w=5.3e-05 

m176 3 61 60 3 penh l=2e-06 w=4.9e-05 

m177 61 62 3 3 penh l=2e-06 w=2.3e-05 

m178 3 60 59 3 penh l=2e-06 w=4.8e-05 

m179 59 60 3 3 penh l=2e-06 w=4.8e-05 

m180 3 62 63 3 penh l=2e-06 w=2.2e-05 

m181 64 65 3 3 penh l=2e-06 w=5e-05 

m182 3 63 65 3 penh l=2e-06 w=4.7e-05 

m183 64 65 3 3 penh l=2e-06 w=4.8e-05 

m184 3 65 64 3 penh l=2e-06 w=4.8e-05 

m185 0 64 58 0 nenh l=2e-06 w=4.6e-05 

m186 58 64 0 0 nenh l=2e-06 w=4.8e-05 

m187 0 64 58 0 nenh l=2e-06 w=4.6e-05 

m188 58 64 0 0 nenh l=2e-06 w=4.8e-05 

m189 0 64 58 0 nenh l=2e-06 w=4.8e-05 

m190 58 64 0 0 nenh l=2e-06 w=4.8e-05 

m191 0 64 58 0 nenh l=2e-06 w=4.8e-05 

m192 58 64 0 0 nenh l=2e-06 w=4.6e-05 

m193 0 65 64 0 nenh l=2e-06 w=6e-05 

m194 64 65 0 0 nenh l=2e-06 w=6e-05 

m195 65 63 0 0 nenh l=2e-06 w=5e-05 

m196 0 60 59 0 nenh l=2e-06 w=3.5e-05 

m197 59 60 0 0 nenh l=2e-06 w=3.4e-05 

m198 0 62 63 0 nenh l=2e-06 w=2.4e-05 

m199 0 60 59 0 nenh l=2e-06 w=2.5e-05 

m200 59 60 0 0 nenh l=2e-06 w=2.5e-05 

m201 0 61 60 0 nenh l=2e-06 w=1.6e-05 

m202 61 62 0 0 nenh l=2e-06 w=2.3e-05 

m203 3 67 66 3 penh l=2e-06 w=9.7e-05 

m204 66 67 3 3 penh l=2e-06 w=9.5e-05 

m205 3 67 66 3 penh l=2e-06 w=9.5e-05 

m206 66 67 3 3 penh l=2e-06 w=9.6e-05 

m207 3 67 66 3 penh l=2e-06 w=9.6e-05 

m208 66 67 3 3 penh l=2e-06 w=9.5e-05 

m209 3 67 66 3 penh l=2e-06 w=9.5e-05 

m210 66 67 3 3 penh l=2e-06 w=9.6e-05 

m211 3 68 67 3 penh l=2e-06 w=5.3e-05 

m212 67 68 3 3 penh l=2e-06 w=5.3e-05 

m213 3 69 68 3 penh l=2e-06 w=4.9e-05 

m214 69 70 3 3 penh l=2e-06 w=2.3e-05 

m215 3 68 67 3 penh l=2e-06 w=4.8e-05 

m216 67 68 3 3 penh l=2e-06 w=4.8e-05 

m217 3 70 71 3 penh l=2e-06 w=2.2e-05 

m218 72 73 3 3 penh l=2e-06 w=5e-05 

m219 3 71 73 3 penh l=2e-06 w=4.7e-05 

m220 72 73 3 3 penh l=2e-06 w=4.8e-05 

m221 3 73 72 3 penh l=2e-06 w=4.8e-05 

m222 0 72 66 0 nenh l=2e-06 w=4.6e-05 

m223 66 72 0 0 nenh l=2e-06 w=4.8e-05 

m224 0 72 66 0 nenh l=2e-06 w=4.6e-05 

m225 66 72 0 0 nenh l=2e-06 w=4.8e-05 

m226 0 72 66 0 nenh l=2e-06 w=4.8e-05 

m227 66 72 0 0 nenh l=2e-06 w=4.8e-05 

m228 0 72 66 0 nenh l=2e-06 w=4.8e-05 

m229 66 72 0 0 nenh l=2e-06 w=4.6e-05 

m230 0 73 72 0 nenh l=2e-06 w=6e-05 

m231 72 73 0 0 nenh l=2e-06 w=6e-05 

m232 73 71 0 0 nenh l=2e-06 w=5e-05 

m233 0 68 67 0 nenh l=2e-06 w=3.5e-05 

m234 67 68 0 0 nenh l=2e-06 w=3.4e-05 

m235 0 70 71 0 nenh l=2e-06 w=2.4e-05 

m236 0 68 67 0 nenh l=2e-06 w=2.5e-05 

m237 67 68 0 0 nenh l=2e-06 w=2.5e-05 

m238 0 69 68 0 nenh l=2e-06 w=1.6e-05 

m239 69 70 0 0 nenh l=2e-06 w=2.3e-05 

m240 0 34 74 0 nenh l=2e-06 w=2.9e-05 

m241 74 34 0 0 nenh l=2e-06 w=1.7e-05 

m242 0 34 74 0 nenh l=2e-06 w=2.9e-05 

m243 74 34 0 0 nenh l=2e-06 w=1.7e-05 

m244 0 34 74 0 nenh l=2e-06 w=1.2e-05 

m245 0 34 74 0 nenh l=2e-06 w=1.2e-05 

m246 74 34 3 3 penh l=2e-06 w=2.2e-05 

m247 3 34 74 3 penh l=2e-06 w=3.4e-05 

m248 74 34 3 3 penh l=2e-06 w=2.3e-05 

m249 74 34 3 3 penh l=2e-06 w=2.2e-05 

m250 3 34 74 3 penh l=2e-06 w=3.4e-05 

m251 74 34 3 3 penh l=2e-06 w=2.3e-05 

m252 74 34 3 3 penh l=2e-06 w=2.7e-05 

m253 74 34 3 3 penh l=2e-06 w=2.7e-05 

m254 75 77 76 3 penh l=2e-06 w=6e-06 

m255 76 79 78 3 penh l=2e-06 w=6e-06 

m256 76 81 80 3 penh l=2e-06 w=6e-06 

m257 80 83 82 3 penh l=2e-06 w=6e-06 

m258 82 84 3 3 penh l=2e-06 w=6e-06 

m259 3 80 84 3 penh l=2e-06 w=6e-06 

m260 84 74 3 3 penh l=2e-06 w=6e-06 

m261 3 84 78 3 penh l=2e-06 w=6e-06 

m262 3 78 85 3 penh l=2e-06 w=2.4e-05 

m263 75 79 76 0 nenh l=2e-06 w=4e-06 

m264 76 77 78 0 nenh l=2e-06 w=4e-06 

m265 3 85 86 3 penh l=2e-06 w=2.8e-05 

m266 86 85 3 3 penh l=2e-06 w=3e-05 

m267 86 85 3 3 penh l=2e-06 w=1.8e-05 

m268 76 83 80 0 nenh l=2e-06 w=4e-06 

m269 80 81 87 0 nenh l=2e-06 w=4e-06 

m270 87 84 0 0 nenh l=2e-06 w=4e-06 

m271 0 80 88 0 nenh l=2e-06 w=8e-06 

m272 88 74 84 0 nenh l=2e-06 w=8e-06 

m273 3 85 86 3 penh l=2e-06 w=1.8e-05 

m274 78 84 0 0 nenh l=2e-06 w=4e-06 

m275 0 78 85 0 nenh l=2e-06 w=1.6e-05 

m276 86 85 0 0 nenh l=2e-06 w=1.4e-05 

m277 0 85 86 0 nenh l=2e-06 w=3.1e-05 

m278 86 85 0 0 nenh l=2e-06 w=1.9e-05 

m279 0 90 89 0 nenh l=2e-06 w=1.6e-05 

m280 0 89 91 0 nenh l=2e-06 w=3.1e-05 

m281 92 79 93 0 nenh l=2e-06 w=4e-06 

m282 93 77 90 0 nenh l=2e-06 w=4e-06 

m283 93 83 94 0 nenh l=2e-06 w=4e-06 

m284 94 81 95 0 nenh l=2e-06 w=4e-06 

m285 95 96 0 0 nenh l=2e-06 w=4e-06 

m286 0 94 97 0 nenh l=2e-06 w=8e-06 

m287 97 74 96 0 nenh l=2e-06 w=8e-06 

m288 90 96 0 0 nenh l=2e-06 w=4e-06 

m289 0 89 91 0 nenh l=2e-06 w=1.4e-05 

m290 91 89 0 0 nenh l=2e-06 w=1.9e-05 

m291 92 77 93 3 penh l=2e-06 w=6e-06 

m292 93 79 90 3 penh l=2e-06 w=6e-06 

m293 93 81 94 3 penh l=2e-06 w=6e-06 

m294 94 83 98 3 penh l=2e-06 w=6e-06 

m295 98 96 3 3 penh l=2e-06 w=6e-06 

m296 3 94 96 3 penh l=2e-06 w=6e-06 

m297 96 74 3 3 penh l=2e-06 w=6e-06 

m298 3 96 90 3 penh l=2e-06 w=6e-06 

m299 3 90 89 3 penh l=2e-06 w=2.4e-05 

m300 3 89 91 3 penh l=2e-06 w=1.8e-05 

m301 91 89 3 3 penh l=2e-06 w=3e-05 

m302 3 89 91 3 penh l=2e-06 w=1.8e-05 

m303 91 89 3 3 penh l=2e-06 w=2.8e-05 

m304 99 77 100 3 penh l=2e-06 w=6e-06 

m305 100 79 101 3 penh l=2e-06 w=6e-06 

m306 100 81 102 3 penh l=2e-06 w=6e-06 

m307 102 83 103 3 penh l=2e-06 w=6e-06 

m308 103 104 3 3 penh l=2e-06 w=6e-06 

m309 3 102 104 3 penh l=2e-06 w=6e-06 

m310 104 74 3 3 penh l=2e-06 w=6e-06 

m311 3 104 101 3 penh l=2e-06 w=6e-06 

m312 3 101 105 3 penh l=2e-06 w=2.4e-05 

m313 99 79 100 0 nenh l=2e-06 w=4e-06 

m314 100 77 101 0 nenh l=2e-06 w=4e-06 

m315 3 105 106 3 penh l=2e-06 w=2.8e-05 

m316 106 105 3 3 penh l=2e-06 w=3e-05 

m317 106 105 3 3 penh l=2e-06 w=1.8e-05 

m318 100 83 102 0 nenh l=2e-06 w=4e-06 

m319 102 81 107 0 nenh l=2e-06 w=4e-06 

m320 107 104 0 0 nenh l=2e-06 w=4e-06 

m321 0 102 108 0 nenh l=2e-06 w=8e-06 

m322 108 74 104 0 nenh l=2e-06 w=8e-06 

m323 3 105 106 3 penh l=2e-06 w=1.8e-05 

m324 101 104 0 0 nenh l=2e-06 w=4e-06 

m325 0 101 105 0 nenh l=2e-06 w=1.6e-05 

m326 106 105 0 0 nenh l=2e-06 w=1.4e-05 

m327 0 105 106 0 nenh l=2e-06 w=3.1e-05 

m328 106 105 0 0 nenh l=2e-06 w=1.9e-05 

m329 0 110 109 0 nenh l=2e-06 w=1.6e-05 

m330 0 109 111 0 nenh l=2e-06 w=3.1e-05 

m331 112 79 113 0 nenh l=2e-06 w=4e-06 

m332 113 77 110 0 nenh l=2e-06 w=4e-06 

m333 113 83 114 0 nenh l=2e-06 w=4e-06 

m334 114 81 115 0 nenh l=2e-06 w=4e-06 

m335 115 116 0 0 nenh l=2e-06 w=4e-06 

m336 0 114 117 0 nenh l=2e-06 w=8e-06 

m337 117 74 116 0 nenh l=2e-06 w=8e-06 

m338 110 116 0 0 nenh l=2e-06 w=4e-06 

m339 0 109 111 0 nenh l=2e-06 w=1.4e-05 

m340 111 109 0 0 nenh l=2e-06 w=1.9e-05 

m341 112 77 113 3 penh l=2e-06 w=6e-06 

m342 113 79 110 3 penh l=2e-06 w=6e-06 

m343 113 81 114 3 penh l=2e-06 w=6e-06 

m344 114 83 118 3 penh l=2e-06 w=6e-06 

m345 118 116 3 3 penh l=2e-06 w=6e-06 

m346 3 114 116 3 penh l=2e-06 w=6e-06 

m347 116 74 3 3 penh l=2e-06 w=6e-06 

m348 3 116 110 3 penh l=2e-06 w=6e-06 

m349 3 110 109 3 penh l=2e-06 w=2.4e-05 

m350 3 109 111 3 penh l=2e-06 w=1.8e-05 

m351 111 109 3 3 penh l=2e-06 w=3e-05 

m352 3 109 111 3 penh l=2e-06 w=1.8e-05 

m353 111 109 3 3 penh l=2e-06 w=2.8e-05 

m354 119 77 120 3 penh l=2e-06 w=6e-06 

m355 120 79 121 3 penh l=2e-06 w=6e-06 

m356 120 81 122 3 penh l=2e-06 w=6e-06 

m357 122 83 123 3 penh l=2e-06 w=6e-06 

m358 123 124 3 3 penh l=2e-06 w=6e-06 

m359 3 122 124 3 penh l=2e-06 w=6e-06 

m360 124 74 3 3 penh l=2e-06 w=6e-06 

m361 3 124 121 3 penh l=2e-06 w=6e-06 

m362 3 121 125 3 penh l=2e-06 w=2.4e-05 

m363 119 79 120 0 nenh l=2e-06 w=4e-06 

m364 120 77 121 0 nenh l=2e-06 w=4e-06 

m365 3 125 126 3 penh l=2e-06 w=2.8e-05 

m366 126 125 3 3 penh l=2e-06 w=3e-05 

m367 126 125 3 3 penh l=2e-06 w=1.8e-05 

m368 120 83 122 0 nenh l=2e-06 w=4e-06 

m369 122 81 127 0 nenh l=2e-06 w=4e-06 

m370 127 124 0 0 nenh l=2e-06 w=4e-06 

m371 0 122 128 0 nenh l=2e-06 w=8e-06 

m372 128 74 124 0 nenh l=2e-06 w=8e-06 

m373 3 125 126 3 penh l=2e-06 w=1.8e-05 

m374 121 124 0 0 nenh l=2e-06 w=4e-06 

m375 0 121 125 0 nenh l=2e-06 w=1.6e-05 

m376 126 125 0 0 nenh l=2e-06 w=1.4e-05 

m377 0 125 126 0 nenh l=2e-06 w=3.1e-05 

m378 126 125 0 0 nenh l=2e-06 w=1.9e-05 

m379 0 130 129 0 nenh l=2e-06 w=1.6e-05 

m380 0 129 131 0 nenh l=2e-06 w=3.1e-05 

m381 132 79 133 0 nenh l=2e-06 w=4e-06 

m382 133 77 130 0 nenh l=2e-06 w=4e-06 

m383 133 83 134 0 nenh l=2e-06 w=4e-06 

m384 134 81 135 0 nenh l=2e-06 w=4e-06 

m385 135 136 0 0 nenh l=2e-06 w=4e-06 

m386 0 134 137 0 nenh l=2e-06 w=8e-06 

m387 137 74 136 0 nenh l=2e-06 w=8e-06 

m388 130 136 0 0 nenh l=2e-06 w=4e-06 

m389 0 129 131 0 nenh l=2e-06 w=1.4e-05 

m390 131 129 0 0 nenh l=2e-06 w=1.9e-05 

m391 132 77 133 3 penh l=2e-06 w=6e-06 

m392 133 79 130 3 penh l=2e-06 w=6e-06 

m393 133 81 134 3 penh l=2e-06 w=6e-06 

m394 134 83 138 3 penh l=2e-06 w=6e-06 

m395 138 136 3 3 penh l=2e-06 w=6e-06 

m396 3 134 136 3 penh l=2e-06 w=6e-06 

m397 136 74 3 3 penh l=2e-06 w=6e-06 

m398 3 136 130 3 penh l=2e-06 w=6e-06 

m399 3 130 129 3 penh l=2e-06 w=2.4e-05 

m400 3 129 131 3 penh l=2e-06 w=1.8e-05 

m401 131 129 3 3 penh l=2e-06 w=3e-05 

m402 3 129 131 3 penh l=2e-06 w=1.8e-05 

m403 131 129 3 3 penh l=2e-06 w=2.8e-05 

m404 139 77 140 3 penh l=2e-06 w=6e-06 

m405 140 79 141 3 penh l=2e-06 w=6e-06 

m406 140 81 142 3 penh l=2e-06 w=6e-06 

m407 142 83 143 3 penh l=2e-06 w=6e-06 

m408 143 144 3 3 penh l=2e-06 w=6e-06 

m409 3 142 144 3 penh l=2e-06 w=6e-06 

m410 144 74 3 3 penh l=2e-06 w=6e-06 

m411 3 144 141 3 penh l=2e-06 w=6e-06 

m412 3 141 145 3 penh l=2e-06 w=2.4e-05 

m413 139 79 140 0 nenh l=2e-06 w=4e-06 

m414 140 77 141 0 nenh l=2e-06 w=4e-06 

m415 3 145 146 3 penh l=2e-06 w=2.8e-05 

m416 146 145 3 3 penh l=2e-06 w=3e-05 

m417 146 145 3 3 penh l=2e-06 w=1.8e-05 

m418 140 83 142 0 nenh l=2e-06 w=4e-06 

m419 142 81 147 0 nenh l=2e-06 w=4e-06 

m420 147 144 0 0 nenh l=2e-06 w=4e-06 

m421 0 142 148 0 nenh l=2e-06 w=8e-06 

m422 148 74 144 0 nenh l=2e-06 w=8e-06 

m423 3 145 146 3 penh l=2e-06 w=1.8e-05 

m424 141 144 0 0 nenh l=2e-06 w=4e-06 

m425 0 141 145 0 nenh l=2e-06 w=1.6e-05 

m426 146 145 0 0 nenh l=2e-06 w=1.4e-05 

m427 0 145 146 0 nenh l=2e-06 w=3.1e-05 

m428 146 145 0 0 nenh l=2e-06 w=1.9e-05 

m429 0 150 149 0 nenh l=2e-06 w=1.6e-05 

m430 0 149 151 0 nenh l=2e-06 w=3.1e-05 

m431 152 79 153 0 nenh l=2e-06 w=4e-06 

m432 153 77 150 0 nenh l=2e-06 w=4e-06 

m433 153 83 154 0 nenh l=2e-06 w=4e-06 

m434 154 81 155 0 nenh l=2e-06 w=4e-06 

m435 155 156 0 0 nenh l=2e-06 w=4e-06 

m436 0 154 157 0 nenh l=2e-06 w=8e-06 

m437 157 74 156 0 nenh l=2e-06 w=8e-06 

m438 150 156 0 0 nenh l=2e-06 w=4e-06 

m439 0 149 151 0 nenh l=2e-06 w=1.4e-05 

m440 151 149 0 0 nenh l=2e-06 w=1.9e-05 

m441 152 77 153 3 penh l=2e-06 w=6e-06 

m442 153 79 150 3 penh l=2e-06 w=6e-06 

m443 153 81 154 3 penh l=2e-06 w=6e-06 

m444 154 83 158 3 penh l=2e-06 w=6e-06 

m445 158 156 3 3 penh l=2e-06 w=6e-06 

m446 3 154 156 3 penh l=2e-06 w=6e-06 

m447 156 74 3 3 penh l=2e-06 w=6e-06 

m448 3 156 150 3 penh l=2e-06 w=6e-06 

m449 3 150 149 3 penh l=2e-06 w=2.4e-05 

m450 3 149 151 3 penh l=2e-06 w=1.8e-05 

m451 151 149 3 3 penh l=2e-06 w=3e-05 

m452 3 149 151 3 penh l=2e-06 w=1.8e-05 

m453 151 149 3 3 penh l=2e-06 w=2.8e-05 

m454 159 77 160 3 penh l=2e-06 w=6e-06 

m455 160 79 161 3 penh l=2e-06 w=6e-06 

m456 160 81 162 3 penh l=2e-06 w=6e-06 

m457 162 83 163 3 penh l=2e-06 w=6e-06 

m458 163 164 3 3 penh l=2e-06 w=6e-06 

m459 3 162 164 3 penh l=2e-06 w=6e-06 

m460 164 74 3 3 penh l=2e-06 w=6e-06 

m461 3 164 161 3 penh l=2e-06 w=6e-06 

m462 3 161 165 3 penh l=2e-06 w=2.4e-05 

m463 159 79 160 0 nenh l=2e-06 w=4e-06 

m464 160 77 161 0 nenh l=2e-06 w=4e-06 

m465 3 165 166 3 penh l=2e-06 w=2.8e-05 

m466 166 165 3 3 penh l=2e-06 w=3e-05 

m467 166 165 3 3 penh l=2e-06 w=1.8e-05 

m468 160 83 162 0 nenh l=2e-06 w=4e-06 

m469 162 81 167 0 nenh l=2e-06 w=4e-06 

m470 167 164 0 0 nenh l=2e-06 w=4e-06 

m471 0 162 168 0 nenh l=2e-06 w=8e-06 

m472 168 74 164 0 nenh l=2e-06 w=8e-06 

m473 3 165 166 3 penh l=2e-06 w=1.8e-05 

m474 161 164 0 0 nenh l=2e-06 w=4e-06 

m475 0 161 165 0 nenh l=2e-06 w=1.6e-05 

m476 166 165 0 0 nenh l=2e-06 w=1.4e-05 

m477 0 165 166 0 nenh l=2e-06 w=3.1e-05 

m478 166 165 0 0 nenh l=2e-06 w=1.9e-05 

m479 0 170 169 0 nenh l=2e-06 w=1.6e-05 

m480 0 169 171 0 nenh l=2e-06 w=3.1e-05 

m481 53 79 172 0 nenh l=2e-06 w=4e-06 

m482 172 77 170 0 nenh l=2e-06 w=4e-06 

m483 172 83 173 0 nenh l=2e-06 w=4e-06 

m484 173 81 174 0 nenh l=2e-06 w=4e-06 

m485 174 175 0 0 nenh l=2e-06 w=4e-06 

m486 0 173 176 0 nenh l=2e-06 w=8e-06 

m487 176 74 175 0 nenh l=2e-06 w=8e-06 

m488 170 175 0 0 nenh l=2e-06 w=4e-06 

m489 0 169 171 0 nenh l=2e-06 w=1.4e-05 

m490 171 169 0 0 nenh l=2e-06 w=1.9e-05 

m491 53 77 172 3 penh l=2e-06 w=6e-06 

m492 172 79 170 3 penh l=2e-06 w=6e-06 

m493 172 81 173 3 penh l=2e-06 w=6e-06 

m494 173 83 177 3 penh l=2e-06 w=6e-06 

m495 177 175 3 3 penh l=2e-06 w=6e-06 

m496 3 173 175 3 penh l=2e-06 w=6e-06 

m497 175 74 3 3 penh l=2e-06 w=6e-06 

m498 3 175 170 3 penh l=2e-06 w=6e-06 

m499 3 170 169 3 penh l=2e-06 w=2.4e-05 

m500 3 169 171 3 penh l=2e-06 w=1.8e-05 

m501 171 169 3 3 penh l=2e-06 w=3e-05 

m502 3 169 171 3 penh l=2e-06 w=1.8e-05 

m503 171 169 3 3 penh l=2e-06 w=2.8e-05 

m504 178 77 179 3 penh l=2e-06 w=6e-06 

m505 179 79 180 3 penh l=2e-06 w=6e-06 

m506 179 81 181 3 penh l=2e-06 w=6e-06 

m507 181 83 182 3 penh l=2e-06 w=6e-06 

m508 182 183 3 3 penh l=2e-06 w=6e-06 

m509 3 181 183 3 penh l=2e-06 w=6e-06 

m510 183 74 3 3 penh l=2e-06 w=6e-06 

m511 3 183 180 3 penh l=2e-06 w=6e-06 

m512 3 180 184 3 penh l=2e-06 w=2.4e-05 

m513 178 79 179 0 nenh l=2e-06 w=4e-06 

m514 179 77 180 0 nenh l=2e-06 w=4e-06 

m515 3 184 185 3 penh l=2e-06 w=2.8e-05 

m516 185 184 3 3 penh l=2e-06 w=3e-05 

m517 185 184 3 3 penh l=2e-06 w=1.8e-05 

m518 179 83 181 0 nenh l=2e-06 w=4e-06 

m519 181 81 186 0 nenh l=2e-06 w=4e-06 

m520 186 183 0 0 nenh l=2e-06 w=4e-06 

m521 0 181 187 0 nenh l=2e-06 w=8e-06 

m522 187 74 183 0 nenh l=2e-06 w=8e-06 

m523 3 184 185 3 penh l=2e-06 w=1.8e-05 

m524 180 183 0 0 nenh l=2e-06 w=4e-06 

m525 0 180 184 0 nenh l=2e-06 w=1.6e-05 

m526 185 184 0 0 nenh l=2e-06 w=1.4e-05 

m527 0 184 185 0 nenh l=2e-06 w=3.1e-05 

m528 185 184 0 0 nenh l=2e-06 w=1.9e-05 

m529 0 189 188 0 nenh l=2e-06 w=1.6e-05 

m530 0 188 190 0 nenh l=2e-06 w=3.1e-05 

m531 48 79 191 0 nenh l=2e-06 w=4e-06 

m532 191 77 189 0 nenh l=2e-06 w=4e-06 

m533 191 83 192 0 nenh l=2e-06 w=4e-06 

m534 192 81 193 0 nenh l=2e-06 w=4e-06 

m535 193 194 0 0 nenh l=2e-06 w=4e-06 

m536 0 192 195 0 nenh l=2e-06 w=8e-06 

m537 195 74 194 0 nenh l=2e-06 w=8e-06 

m538 189 194 0 0 nenh l=2e-06 w=4e-06 

m539 0 188 190 0 nenh l=2e-06 w=1.4e-05 

m540 190 188 0 0 nenh l=2e-06 w=1.9e-05 

m541 48 77 191 3 penh l=2e-06 w=6e-06 

m542 191 79 189 3 penh l=2e-06 w=6e-06 

m543 191 81 192 3 penh l=2e-06 w=6e-06 

m544 192 83 196 3 penh l=2e-06 w=6e-06 

m545 196 194 3 3 penh l=2e-06 w=6e-06 

m546 3 192 194 3 penh l=2e-06 w=6e-06 

m547 194 74 3 3 penh l=2e-06 w=6e-06 

m548 3 194 189 3 penh l=2e-06 w=6e-06 

m549 3 189 188 3 penh l=2e-06 w=2.4e-05 

m550 3 188 190 3 penh l=2e-06 w=1.8e-05 

m551 190 188 3 3 penh l=2e-06 w=3e-05 

m552 3 188 190 3 penh l=2e-06 w=1.8e-05 

m553 190 188 3 3 penh l=2e-06 w=2.8e-05 

m554 197 77 198 3 penh l=2e-06 w=6e-06 

m555 198 79 199 3 penh l=2e-06 w=6e-06 

m556 198 81 200 3 penh l=2e-06 w=6e-06 

m557 200 83 201 3 penh l=2e-06 w=6e-06 

m558 201 202 3 3 penh l=2e-06 w=6e-06 

m559 3 200 202 3 penh l=2e-06 w=6e-06 

m560 202 74 3 3 penh l=2e-06 w=6e-06 

m561 3 202 199 3 penh l=2e-06 w=6e-06 

m562 3 199 203 3 penh l=2e-06 w=2.4e-05 

m563 197 79 198 0 nenh l=2e-06 w=4e-06 

m564 198 77 199 0 nenh l=2e-06 w=4e-06 

m565 3 203 204 3 penh l=2e-06 w=2.8e-05 

m566 204 203 3 3 penh l=2e-06 w=3e-05 

m567 204 203 3 3 penh l=2e-06 w=1.8e-05 

m568 198 83 200 0 nenh l=2e-06 w=4e-06 

m569 200 81 205 0 nenh l=2e-06 w=4e-06 

m570 205 202 0 0 nenh l=2e-06 w=4e-06 

m571 0 200 206 0 nenh l=2e-06 w=8e-06 

m572 206 74 202 0 nenh l=2e-06 w=8e-06 

m573 3 203 204 3 penh l=2e-06 w=1.8e-05 

m574 199 202 0 0 nenh l=2e-06 w=4e-06 

m575 0 199 203 0 nenh l=2e-06 w=1.6e-05 

m576 204 203 0 0 nenh l=2e-06 w=1.4e-05 

m577 0 203 204 0 nenh l=2e-06 w=3.1e-05 

m578 204 203 0 0 nenh l=2e-06 w=1.9e-05 

m579 0 208 207 0 nenh l=2e-06 w=1.6e-05 

m580 0 207 209 0 nenh l=2e-06 w=3.1e-05 

m581 43 79 210 0 nenh l=2e-06 w=4e-06 

m582 210 77 208 0 nenh l=2e-06 w=4e-06 

m583 210 83 211 0 nenh l=2e-06 w=4e-06 

m584 211 81 212 0 nenh l=2e-06 w=4e-06 

m585 212 213 0 0 nenh l=2e-06 w=4e-06 

m586 0 211 214 0 nenh l=2e-06 w=8e-06 

m587 214 74 213 0 nenh l=2e-06 w=8e-06 

m588 208 213 0 0 nenh l=2e-06 w=4e-06 

m589 0 207 209 0 nenh l=2e-06 w=1.4e-05 

m590 209 207 0 0 nenh l=2e-06 w=1.9e-05 

m591 43 77 210 3 penh l=2e-06 w=6e-06 

m592 210 79 208 3 penh l=2e-06 w=6e-06 

m593 210 81 211 3 penh l=2e-06 w=6e-06 

m594 211 83 215 3 penh l=2e-06 w=6e-06 

m595 215 213 3 3 penh l=2e-06 w=6e-06 

m596 3 211 213 3 penh l=2e-06 w=6e-06 

m597 213 74 3 3 penh l=2e-06 w=6e-06 

m598 3 213 208 3 penh l=2e-06 w=6e-06 

m599 3 208 207 3 penh l=2e-06 w=2.4e-05 

m600 3 207 209 3 penh l=2e-06 w=1.8e-05 

m601 209 207 3 3 penh l=2e-06 w=3e-05 

m602 3 207 209 3 penh l=2e-06 w=1.8e-05 

m603 209 207 3 3 penh l=2e-06 w=2.8e-05 

m604 216 77 217 3 penh l=2e-06 w=6e-06 

m605 217 79 218 3 penh l=2e-06 w=6e-06 

m606 217 81 219 3 penh l=2e-06 w=6e-06 

m607 219 83 220 3 penh l=2e-06 w=6e-06 

m608 220 221 3 3 penh l=2e-06 w=6e-06 

m609 3 219 221 3 penh l=2e-06 w=6e-06 

m610 221 74 3 3 penh l=2e-06 w=6e-06 

m611 3 221 218 3 penh l=2e-06 w=6e-06 

m612 3 218 222 3 penh l=2e-06 w=2.4e-05 

m613 216 79 217 0 nenh l=2e-06 w=4e-06 

m614 217 77 218 0 nenh l=2e-06 w=4e-06 

m615 3 222 223 3 penh l=2e-06 w=2.8e-05 

m616 223 222 3 3 penh l=2e-06 w=3e-05 

m617 223 222 3 3 penh l=2e-06 w=1.8e-05 

m618 217 83 219 0 nenh l=2e-06 w=4e-06 

m619 219 81 224 0 nenh l=2e-06 w=4e-06 

m620 224 221 0 0 nenh l=2e-06 w=4e-06 

m621 0 219 225 0 nenh l=2e-06 w=8e-06 

m622 225 74 221 0 nenh l=2e-06 w=8e-06 

m623 3 222 223 3 penh l=2e-06 w=1.8e-05 

m624 218 221 0 0 nenh l=2e-06 w=4e-06 

m625 0 218 222 0 nenh l=2e-06 w=1.6e-05 

m626 223 222 0 0 nenh l=2e-06 w=1.4e-05 

m627 0 222 223 0 nenh l=2e-06 w=3.1e-05 

m628 223 222 0 0 nenh l=2e-06 w=1.9e-05 

m629 0 227 226 0 nenh l=2e-06 w=1.6e-05 

m630 0 226 228 0 nenh l=2e-06 w=3.1e-05 

m631 38 79 229 0 nenh l=2e-06 w=4e-06 

m632 229 77 227 0 nenh l=2e-06 w=4e-06 

m633 229 83 230 0 nenh l=2e-06 w=4e-06 

m634 230 81 231 0 nenh l=2e-06 w=4e-06 

m635 231 232 0 0 nenh l=2e-06 w=4e-06 

m636 0 230 233 0 nenh l=2e-06 w=8e-06 

m637 233 74 232 0 nenh l=2e-06 w=8e-06 

m638 227 232 0 0 nenh l=2e-06 w=4e-06 

m639 0 226 228 0 nenh l=2e-06 w=1.4e-05 

m640 228 226 0 0 nenh l=2e-06 w=1.9e-05 

m641 38 77 229 3 penh l=2e-06 w=6e-06 

m642 229 79 227 3 penh l=2e-06 w=6e-06 

m643 229 81 230 3 penh l=2e-06 w=6e-06 

m644 230 83 234 3 penh l=2e-06 w=6e-06 

m645 234 232 3 3 penh l=2e-06 w=6e-06 

m646 3 230 232 3 penh l=2e-06 w=6e-06 

m647 232 74 3 3 penh l=2e-06 w=6e-06 

m648 3 232 227 3 penh l=2e-06 w=6e-06 

m649 3 227 226 3 penh l=2e-06 w=2.4e-05 

m650 3 226 228 3 penh l=2e-06 w=1.8e-05 

m651 228 226 3 3 penh l=2e-06 w=3e-05 

m652 3 226 228 3 penh l=2e-06 w=1.8e-05 

m653 228 226 3 3 penh l=2e-06 w=2.8e-05 

m654 152 235 3 3 penh l=2e-06 w=6.2e-05 

m655 3 236 235 3 penh l=2e-06 w=6.2e-05 

m656 236 237 3 3 penh l=2e-06 w=2.9e-05 

m657 3 238 237 3 penh l=4e-06 w=2.9e-05 

m658 236 237 0 0 nenh l=2e-06 w=2.1e-05 

m659 0 238 237 0 nenh l=4e-06 w=2.1e-05 

m660 152 235 0 0 nenh l=2e-06 w=4.8e-05 

m661 0 236 235 0 nenh l=2e-06 w=4.8e-05 

m662 238 0 0 0 nenh l=4e-06 w=2.5e-05 

m663 3 240 239 3 penh l=2e-06 w=9.7e-05 

m664 239 240 3 3 penh l=2e-06 w=9.5e-05 

m665 3 240 239 3 penh l=2e-06 w=9.5e-05 

m666 239 240 3 3 penh l=2e-06 w=9.6e-05 

m667 3 240 239 3 penh l=2e-06 w=9.6e-05 

m668 239 240 3 3 penh l=2e-06 w=9.5e-05 

m669 3 240 239 3 penh l=2e-06 w=9.5e-05 

m670 239 240 3 3 penh l=2e-06 w=9.6e-05 

m671 3 241 240 3 penh l=2e-06 w=5.3e-05 

m672 240 241 3 3 penh l=2e-06 w=5.3e-05 

m673 3 242 241 3 penh l=2e-06 w=4.9e-05 

m674 242 243 3 3 penh l=2e-06 w=2.3e-05 

m675 3 241 240 3 penh l=2e-06 w=4.8e-05 

m676 240 241 3 3 penh l=2e-06 w=4.8e-05 

m677 3 243 244 3 penh l=2e-06 w=2.2e-05 

m678 245 246 3 3 penh l=2e-06 w=5e-05 

m679 3 244 246 3 penh l=2e-06 w=4.7e-05 

m680 245 246 3 3 penh l=2e-06 w=4.8e-05 

m681 3 246 245 3 penh l=2e-06 w=4.8e-05 

m682 0 245 239 0 nenh l=2e-06 w=4.6e-05 

m683 239 245 0 0 nenh l=2e-06 w=4.8e-05 

m684 0 245 239 0 nenh l=2e-06 w=4.6e-05 

m685 239 245 0 0 nenh l=2e-06 w=4.8e-05 

m686 0 245 239 0 nenh l=2e-06 w=4.8e-05 

m687 239 245 0 0 nenh l=2e-06 w=4.8e-05 

m688 0 245 239 0 nenh l=2e-06 w=4.8e-05 

m689 239 245 0 0 nenh l=2e-06 w=4.6e-05 

m690 0 246 245 0 nenh l=2e-06 w=6e-05 

m691 245 246 0 0 nenh l=2e-06 w=6e-05 

m692 246 244 0 0 nenh l=2e-06 w=5e-05 

m693 0 241 240 0 nenh l=2e-06 w=3.5e-05 

m694 240 241 0 0 nenh l=2e-06 w=3.4e-05 

m695 0 243 244 0 nenh l=2e-06 w=2.4e-05 

m696 0 241 240 0 nenh l=2e-06 w=2.5e-05 

m697 240 241 0 0 nenh l=2e-06 w=2.5e-05 

m698 0 242 241 0 nenh l=2e-06 w=1.6e-05 

m699 242 243 0 0 nenh l=2e-06 w=2.3e-05 

m700 3 248 247 3 penh l=2e-06 w=9.7e-05 

m701 247 248 3 3 penh l=2e-06 w=9.5e-05 

m702 3 248 247 3 penh l=2e-06 w=9.5e-05 

m703 247 248 3 3 penh l=2e-06 w=9.6e-05 

m704 3 248 247 3 penh l=2e-06 w=9.6e-05 

m705 247 248 3 3 penh l=2e-06 w=9.5e-05 

m706 3 248 247 3 penh l=2e-06 w=9.5e-05 

m707 247 248 3 3 penh l=2e-06 w=9.6e-05 

m708 3 249 248 3 penh l=2e-06 w=5.3e-05 

m709 248 249 3 3 penh l=2e-06 w=5.3e-05 

m710 3 250 249 3 penh l=2e-06 w=4.9e-05 

m711 250 251 3 3 penh l=2e-06 w=2.3e-05 

m712 3 249 248 3 penh l=2e-06 w=4.8e-05 

m713 248 249 3 3 penh l=2e-06 w=4.8e-05 

m714 3 251 252 3 penh l=2e-06 w=2.2e-05 

m715 253 254 3 3 penh l=2e-06 w=5e-05 

m716 3 252 254 3 penh l=2e-06 w=4.7e-05 

m717 253 254 3 3 penh l=2e-06 w=4.8e-05 

m718 3 254 253 3 penh l=2e-06 w=4.8e-05 

m719 0 253 247 0 nenh l=2e-06 w=4.6e-05 

m720 247 253 0 0 nenh l=2e-06 w=4.8e-05 

m721 0 253 247 0 nenh l=2e-06 w=4.6e-05 

m722 247 253 0 0 nenh l=2e-06 w=4.8e-05 

m723 0 253 247 0 nenh l=2e-06 w=4.8e-05 

m724 247 253 0 0 nenh l=2e-06 w=4.8e-05 

m725 0 253 247 0 nenh l=2e-06 w=4.8e-05 

m726 247 253 0 0 nenh l=2e-06 w=4.6e-05 

m727 0 254 253 0 nenh l=2e-06 w=6e-05 

m728 253 254 0 0 nenh l=2e-06 w=6e-05 

m729 254 252 0 0 nenh l=2e-06 w=5e-05 

m730 0 249 248 0 nenh l=2e-06 w=3.5e-05 

m731 248 249 0 0 nenh l=2e-06 w=3.4e-05 

m732 0 251 252 0 nenh l=2e-06 w=2.4e-05 

m733 0 249 248 0 nenh l=2e-06 w=2.5e-05 

m734 248 249 0 0 nenh l=2e-06 w=2.5e-05 

m735 0 250 249 0 nenh l=2e-06 w=1.6e-05 

m736 250 251 0 0 nenh l=2e-06 w=2.3e-05 

m737 3 256 255 3 penh l=2e-06 w=9.7e-05 

m738 255 256 3 3 penh l=2e-06 w=9.5e-05 

m739 3 256 255 3 penh l=2e-06 w=9.5e-05 

m740 255 256 3 3 penh l=2e-06 w=9.6e-05 

m741 3 256 255 3 penh l=2e-06 w=9.6e-05 

m742 255 256 3 3 penh l=2e-06 w=9.5e-05 

m743 3 256 255 3 penh l=2e-06 w=9.5e-05 

m744 255 256 3 3 penh l=2e-06 w=9.6e-05 

m745 3 257 256 3 penh l=2e-06 w=5.3e-05 

m746 256 257 3 3 penh l=2e-06 w=5.3e-05 

m747 3 258 257 3 penh l=2e-06 w=4.9e-05 

m748 258 259 3 3 penh l=2e-06 w=2.3e-05 

m749 3 257 256 3 penh l=2e-06 w=4.8e-05 

m750 256 257 3 3 penh l=2e-06 w=4.8e-05 

m751 3 259 260 3 penh l=2e-06 w=2.2e-05 

m752 261 262 3 3 penh l=2e-06 w=5e-05 

m753 3 260 262 3 penh l=2e-06 w=4.7e-05 

m754 261 262 3 3 penh l=2e-06 w=4.8e-05 

m755 3 262 261 3 penh l=2e-06 w=4.8e-05 

m756 0 261 255 0 nenh l=2e-06 w=4.6e-05 

m757 255 261 0 0 nenh l=2e-06 w=4.8e-05 

m758 0 261 255 0 nenh l=2e-06 w=4.6e-05 

m759 255 261 0 0 nenh l=2e-06 w=4.8e-05 

m760 0 261 255 0 nenh l=2e-06 w=4.8e-05 

m761 255 261 0 0 nenh l=2e-06 w=4.8e-05 

m762 0 261 255 0 nenh l=2e-06 w=4.8e-05 

m763 255 261 0 0 nenh l=2e-06 w=4.6e-05 

m764 0 262 261 0 nenh l=2e-06 w=6e-05 

m765 261 262 0 0 nenh l=2e-06 w=6e-05 

m766 262 260 0 0 nenh l=2e-06 w=5e-05 

m767 0 257 256 0 nenh l=2e-06 w=3.5e-05 

m768 256 257 0 0 nenh l=2e-06 w=3.4e-05 

m769 0 259 260 0 nenh l=2e-06 w=2.4e-05 

m770 0 257 256 0 nenh l=2e-06 w=2.5e-05 

m771 256 257 0 0 nenh l=2e-06 w=2.5e-05 

m772 0 258 257 0 nenh l=2e-06 w=1.6e-05 

m773 258 259 0 0 nenh l=2e-06 w=2.3e-05 

m774 3 264 263 3 penh l=2e-06 w=9.7e-05 

m775 263 264 3 3 penh l=2e-06 w=9.5e-05 

m776 3 264 263 3 penh l=2e-06 w=9.5e-05 

m777 263 264 3 3 penh l=2e-06 w=9.6e-05 

m778 3 264 263 3 penh l=2e-06 w=9.6e-05 

m779 263 264 3 3 penh l=2e-06 w=9.5e-05 

m780 3 264 263 3 penh l=2e-06 w=9.5e-05 

m781 263 264 3 3 penh l=2e-06 w=9.6e-05 

m782 3 265 264 3 penh l=2e-06 w=5.3e-05 

m783 264 265 3 3 penh l=2e-06 w=5.3e-05 

m784 3 266 265 3 penh l=2e-06 w=4.9e-05 

m785 266 267 3 3 penh l=2e-06 w=2.3e-05 

m786 3 265 264 3 penh l=2e-06 w=4.8e-05 

m787 264 265 3 3 penh l=2e-06 w=4.8e-05 

m788 3 267 268 3 penh l=2e-06 w=2.2e-05 

m789 269 270 3 3 penh l=2e-06 w=5e-05 

m790 3 268 270 3 penh l=2e-06 w=4.7e-05 

m791 269 270 3 3 penh l=2e-06 w=4.8e-05 

m792 3 270 269 3 penh l=2e-06 w=4.8e-05 

m793 0 269 263 0 nenh l=2e-06 w=4.6e-05 

m794 263 269 0 0 nenh l=2e-06 w=4.8e-05 

m795 0 269 263 0 nenh l=2e-06 w=4.6e-05 

m796 263 269 0 0 nenh l=2e-06 w=4.8e-05 

m797 0 269 263 0 nenh l=2e-06 w=4.8e-05 

m798 263 269 0 0 nenh l=2e-06 w=4.8e-05 

m799 0 269 263 0 nenh l=2e-06 w=4.8e-05 

m800 263 269 0 0 nenh l=2e-06 w=4.6e-05 

m801 0 270 269 0 nenh l=2e-06 w=6e-05 

m802 269 270 0 0 nenh l=2e-06 w=6e-05 

m803 270 268 0 0 nenh l=2e-06 w=5e-05 

m804 0 265 264 0 nenh l=2e-06 w=3.5e-05 

m805 264 265 0 0 nenh l=2e-06 w=3.4e-05 

m806 0 267 268 0 nenh l=2e-06 w=2.4e-05 

m807 0 265 264 0 nenh l=2e-06 w=2.5e-05 

m808 264 265 0 0 nenh l=2e-06 w=2.5e-05 

m809 0 266 265 0 nenh l=2e-06 w=1.6e-05 

m810 266 267 0 0 nenh l=2e-06 w=2.3e-05 

m811 271 273 272 0 nenh l=2e-06 w=4e-06 

m812 272 275 274 0 nenh l=2e-06 w=4e-06 

m813 276 272 0 0 nenh l=2e-06 w=4e-06 

m814 0 276 277 0 nenh l=2e-06 w=1.2e-05 

m815 271 275 272 3 penh l=2e-06 w=6e-06 

m816 272 273 274 3 penh l=2e-06 w=6e-06 

m817 276 272 3 3 penh l=2e-06 w=6e-06 

m818 3 276 277 3 penh l=2e-06 w=1.8e-05 

m819 278 273 279 0 nenh l=2e-06 w=4e-06 

m820 279 275 280 0 nenh l=2e-06 w=4e-06 

m821 281 279 0 0 nenh l=2e-06 w=4e-06 

m822 0 281 282 0 nenh l=2e-06 w=1.2e-05 

m823 278 275 279 3 penh l=2e-06 w=6e-06 

m824 279 273 280 3 penh l=2e-06 w=6e-06 

m825 281 279 3 3 penh l=2e-06 w=6e-06 

m826 3 281 282 3 penh l=2e-06 w=1.8e-05 

m827 283 273 284 0 nenh l=2e-06 w=4e-06 

m828 284 275 285 0 nenh l=2e-06 w=4e-06 

m829 286 284 0 0 nenh l=2e-06 w=4e-06 

m830 0 286 287 0 nenh l=2e-06 w=1.2e-05 

m831 283 275 284 3 penh l=2e-06 w=6e-06 

m832 284 273 285 3 penh l=2e-06 w=6e-06 

m833 286 284 3 3 penh l=2e-06 w=6e-06 

m834 3 286 287 3 penh l=2e-06 w=1.8e-05 

m835 288 273 289 0 nenh l=2e-06 w=4e-06 

m836 289 275 290 0 nenh l=2e-06 w=4e-06 

m837 291 289 0 0 nenh l=2e-06 w=4e-06 

m838 0 291 292 0 nenh l=2e-06 w=1.2e-05 

m839 288 275 289 3 penh l=2e-06 w=6e-06 

m840 289 273 290 3 penh l=2e-06 w=6e-06 

m841 291 289 3 3 penh l=2e-06 w=6e-06 

m842 3 291 292 3 penh l=2e-06 w=1.8e-05 

m843 293 273 294 0 nenh l=2e-06 w=4e-06 

m844 294 275 295 0 nenh l=2e-06 w=4e-06 

m845 296 294 0 0 nenh l=2e-06 w=4e-06 

m846 0 296 267 0 nenh l=2e-06 w=1.2e-05 

m847 293 275 294 3 penh l=2e-06 w=6e-06 

m848 294 273 295 3 penh l=2e-06 w=6e-06 

m849 296 294 3 3 penh l=2e-06 w=6e-06 

m850 3 296 267 3 penh l=2e-06 w=1.8e-05 

m851 297 273 298 0 nenh l=2e-06 w=4e-06 

m852 298 275 299 0 nenh l=2e-06 w=4e-06 

m853 300 298 0 0 nenh l=2e-06 w=4e-06 

m854 0 300 259 0 nenh l=2e-06 w=1.2e-05 

m855 297 275 298 3 penh l=2e-06 w=6e-06 

m856 298 273 299 3 penh l=2e-06 w=6e-06 

m857 300 298 3 3 penh l=2e-06 w=6e-06 

m858 3 300 259 3 penh l=2e-06 w=1.8e-05 

m859 301 273 302 0 nenh l=2e-06 w=4e-06 

m860 302 275 303 0 nenh l=2e-06 w=4e-06 

m861 304 302 0 0 nenh l=2e-06 w=4e-06 

m862 0 304 251 0 nenh l=2e-06 w=1.2e-05 

m863 301 275 302 3 penh l=2e-06 w=6e-06 

m864 302 273 303 3 penh l=2e-06 w=6e-06 

m865 304 302 3 3 penh l=2e-06 w=6e-06 

m866 3 304 251 3 penh l=2e-06 w=1.8e-05 

m867 305 273 306 0 nenh l=2e-06 w=4e-06 

m868 306 275 307 0 nenh l=2e-06 w=4e-06 

m869 308 306 0 0 nenh l=2e-06 w=4e-06 

m870 0 308 243 0 nenh l=2e-06 w=1.2e-05 

m871 305 275 306 3 penh l=2e-06 w=6e-06 

m872 306 273 307 3 penh l=2e-06 w=6e-06 

m873 308 306 3 3 penh l=2e-06 w=6e-06 

m874 3 308 243 3 penh l=2e-06 w=1.8e-05 

m875 309 273 310 0 nenh l=2e-06 w=4e-06 

m876 310 275 311 0 nenh l=2e-06 w=4e-06 

m877 312 310 0 0 nenh l=2e-06 w=4e-06 

m878 0 312 70 0 nenh l=2e-06 w=1.2e-05 

m879 309 275 310 3 penh l=2e-06 w=6e-06 

m880 310 273 311 3 penh l=2e-06 w=6e-06 

m881 312 310 3 3 penh l=2e-06 w=6e-06 

m882 3 312 70 3 penh l=2e-06 w=1.8e-05 

m883 313 273 314 0 nenh l=2e-06 w=4e-06 

m884 314 275 315 0 nenh l=2e-06 w=4e-06 

m885 316 314 0 0 nenh l=2e-06 w=4e-06 

m886 0 316 62 0 nenh l=2e-06 w=1.2e-05 

m887 313 275 314 3 penh l=2e-06 w=6e-06 

m888 314 273 315 3 penh l=2e-06 w=6e-06 

m889 316 314 3 3 penh l=2e-06 w=6e-06 

m890 3 316 62 3 penh l=2e-06 w=1.8e-05 

m891 317 273 318 0 nenh l=2e-06 w=4e-06 

m892 318 275 319 0 nenh l=2e-06 w=4e-06 

m893 320 318 0 0 nenh l=2e-06 w=4e-06 

m894 0 320 8 0 nenh l=2e-06 w=1.2e-05 

m895 317 275 318 3 penh l=2e-06 w=6e-06 

m896 318 273 319 3 penh l=2e-06 w=6e-06 

m897 320 318 3 3 penh l=2e-06 w=6e-06 

m898 3 320 8 3 penh l=2e-06 w=1.8e-05 

m899 16 322 321 0 nenh l=2e-06 w=4e-06 

m900 321 16 322 0 nenh l=2e-06 w=4e-06 

m901 322 24 0 0 nenh l=2e-06 w=4e-06 

m902 0 321 323 0 nenh l=2e-06 w=4e-06 

m903 324 323 0 0 nenh l=2e-06 w=4e-06 

m904 0 324 275 0 nenh l=2e-06 w=1.2e-05 

m905 0 323 273 0 nenh l=2e-06 w=1.2e-05 

m906 16 24 321 3 penh l=2e-06 w=6e-06 

m907 321 16 24 3 penh l=2e-06 w=6e-06 

m908 322 24 3 3 penh l=2e-06 w=6e-06 

m909 3 321 323 3 penh l=2e-06 w=6e-06 

m910 324 323 3 3 penh l=2e-06 w=6e-06 

m911 3 324 275 3 penh l=2e-06 w=1.8e-05 

m912 3 323 273 3 penh l=2e-06 w=1.8e-05 

m913 325 327 326 3 penh l=2e-06 w=5e-06 

m914 326 329 328 3 penh l=2e-06 w=5e-06 

m915 328 330 3 3 penh l=2e-06 w=5e-06 

m916 3 326 330 3 penh l=2e-06 w=6e-06 

m917 330 28 3 3 penh l=2e-06 w=6e-06 

m918 3 330 309 3 penh l=2e-06 w=2.5e-05 

m919 325 329 326 0 nenh l=2e-06 w=5e-06 

m920 326 327 331 0 nenh l=2e-06 w=5e-06 

m921 331 330 0 0 nenh l=2e-06 w=5e-06 

m922 0 326 332 0 nenh l=2e-06 w=1.3e-05 

m923 332 28 330 0 nenh l=2e-06 w=1.2e-05 

m924 0 330 309 0 nenh l=2e-06 w=1.4e-05 

m925 333 327 334 3 penh l=2e-06 w=5e-06 

m926 334 329 335 3 penh l=2e-06 w=5e-06 

m927 335 336 3 3 penh l=2e-06 w=5e-06 

m928 3 334 336 3 penh l=2e-06 w=6e-06 

m929 336 28 3 3 penh l=2e-06 w=6e-06 

m930 3 336 313 3 penh l=2e-06 w=2.5e-05 

m931 333 329 334 0 nenh l=2e-06 w=5e-06 

m932 334 327 337 0 nenh l=2e-06 w=5e-06 

m933 337 336 0 0 nenh l=2e-06 w=5e-06 

m934 0 334 338 0 nenh l=2e-06 w=1.3e-05 

m935 338 28 336 0 nenh l=2e-06 w=1.2e-05 

m936 0 336 313 0 nenh l=2e-06 w=1.4e-05 

m937 339 327 340 3 penh l=2e-06 w=5e-06 

m938 340 329 341 3 penh l=2e-06 w=5e-06 

m939 341 342 3 3 penh l=2e-06 w=5e-06 

m940 3 340 342 3 penh l=2e-06 w=6e-06 

m941 342 28 3 3 penh l=2e-06 w=6e-06 

m942 3 342 317 3 penh l=2e-06 w=2.5e-05 

m943 339 329 340 0 nenh l=2e-06 w=5e-06 

m944 340 327 343 0 nenh l=2e-06 w=5e-06 

m945 343 342 0 0 nenh l=2e-06 w=5e-06 

m946 0 340 344 0 nenh l=2e-06 w=1.3e-05 

m947 344 28 342 0 nenh l=2e-06 w=1.2e-05 

m948 0 342 317 0 nenh l=2e-06 w=1.4e-05 

m949 345 327 346 3 penh l=2e-06 w=5e-06 

m950 346 329 347 3 penh l=2e-06 w=5e-06 

m951 347 348 3 3 penh l=2e-06 w=5e-06 

m952 3 346 348 3 penh l=2e-06 w=6e-06 

m953 348 28 3 3 penh l=2e-06 w=6e-06 

m954 3 348 16 3 penh l=2e-06 w=2.5e-05 

m955 345 329 346 0 nenh l=2e-06 w=5e-06 

m956 346 327 349 0 nenh l=2e-06 w=5e-06 

m957 349 348 0 0 nenh l=2e-06 w=5e-06 

m958 0 346 350 0 nenh l=2e-06 w=1.3e-05 

m959 350 28 348 0 nenh l=2e-06 w=1.2e-05 

m960 0 348 16 0 nenh l=2e-06 w=1.4e-05 

m961 351 327 352 3 penh l=2e-06 w=5e-06 

m962 352 329 353 3 penh l=2e-06 w=5e-06 

m963 353 354 3 3 penh l=2e-06 w=5e-06 

m964 3 352 354 3 penh l=2e-06 w=6e-06 

m965 354 28 3 3 penh l=2e-06 w=6e-06 

m966 3 354 24 3 penh l=2e-06 w=2.5e-05 

m967 351 329 352 0 nenh l=2e-06 w=5e-06 

m968 352 327 355 0 nenh l=2e-06 w=5e-06 

m969 355 354 0 0 nenh l=2e-06 w=5e-06 

m970 0 352 356 0 nenh l=2e-06 w=1.3e-05 

m971 356 28 354 0 nenh l=2e-06 w=1.2e-05 

m972 0 354 24 0 nenh l=2e-06 w=1.4e-05 

m973 357 359 358 0 nenh l=2e-06 w=1.2e-05 

m974 357 361 360 0 nenh l=2e-06 w=1.2e-05 

m975 360 363 362 0 nenh l=2e-06 w=1.2e-05 

m976 362 365 364 0 nenh l=2e-06 w=1.4e-05 

m977 0 358 366 0 nenh l=2e-06 w=6e-06 

m978 3 329 358 3 penh l=2e-06 w=1e-05 

m979 358 366 3 3 penh l=8e-06 w=4e-06 

m980 3 358 366 3 penh l=2e-06 w=1.6e-05 

m981 3 368 367 3 penh l=2e-06 w=1.6e-05 

m982 3 329 368 3 penh l=2e-06 w=1e-05 

m983 368 367 3 3 penh l=8e-06 w=4e-06 

m984 367 368 0 0 nenh l=2e-06 w=6e-06 

m985 0 329 364 0 nenh l=2e-06 w=1.4e-05 

m986 369 370 364 0 nenh l=2e-06 w=8e-06 

m987 364 361 371 0 nenh l=2e-06 w=1e-05 

m988 371 373 372 0 nenh l=2e-06 w=1e-05 

m989 372 374 364 0 nenh l=2e-06 w=8e-06 

m990 364 375 368 0 nenh l=2e-06 w=6e-06 

m991 368 365 369 0 nenh l=2e-06 w=6e-06 

m992 369 363 372 0 nenh l=2e-06 w=8e-06 

m993 376 378 377 0 nenh l=2e-06 w=1.2e-05 

m994 376 380 379 0 nenh l=2e-06 w=1.2e-05 

m995 379 382 381 0 nenh l=2e-06 w=1.2e-05 

m996 381 384 383 0 nenh l=2e-06 w=1.4e-05 

m997 0 377 385 0 nenh l=2e-06 w=6e-06 

m998 3 329 377 3 penh l=2e-06 w=1e-05 

m999 377 385 3 3 penh l=8e-06 w=4e-06 

m1000 3 377 385 3 penh l=2e-06 w=1.6e-05 

m1001 3 387 386 3 penh l=2e-06 w=1.6e-05 

m1002 3 329 387 3 penh l=2e-06 w=1e-05 

m1003 387 386 3 3 penh l=8e-06 w=4e-06 

m1004 386 387 0 0 nenh l=2e-06 w=6e-06 

m1005 0 329 383 0 nenh l=2e-06 w=1.4e-05 

m1006 388 389 383 0 nenh l=2e-06 w=8e-06 

m1007 383 380 390 0 nenh l=2e-06 w=1e-05 

m1008 390 392 391 0 nenh l=2e-06 w=1e-05 

m1009 391 393 383 0 nenh l=2e-06 w=8e-06 

m1010 383 394 387 0 nenh l=2e-06 w=6e-06 

m1011 387 384 388 0 nenh l=2e-06 w=6e-06 

m1012 388 382 391 0 nenh l=2e-06 w=8e-06 

m1013 395 397 396 0 nenh l=2e-06 w=1.2e-05 

m1014 395 399 398 0 nenh l=2e-06 w=1.2e-05 

m1015 398 401 400 0 nenh l=2e-06 w=1.2e-05 

m1016 400 403 402 0 nenh l=2e-06 w=1.4e-05 

m1017 0 396 404 0 nenh l=2e-06 w=6e-06 

m1018 3 329 396 3 penh l=2e-06 w=1e-05 

m1019 396 404 3 3 penh l=8e-06 w=4e-06 

m1020 3 396 404 3 penh l=2e-06 w=1.6e-05 

m1021 3 406 405 3 penh l=2e-06 w=1.6e-05 

m1022 3 329 406 3 penh l=2e-06 w=1e-05 

m1023 406 405 3 3 penh l=8e-06 w=4e-06 

m1024 405 406 0 0 nenh l=2e-06 w=6e-06 

m1025 0 329 402 0 nenh l=2e-06 w=1.4e-05 

m1026 407 408 402 0 nenh l=2e-06 w=8e-06 

m1027 402 399 409 0 nenh l=2e-06 w=1e-05 

m1028 409 411 410 0 nenh l=2e-06 w=1e-05 

m1029 410 412 402 0 nenh l=2e-06 w=8e-06 

m1030 402 413 406 0 nenh l=2e-06 w=6e-06 

m1031 406 403 407 0 nenh l=2e-06 w=6e-06 

m1032 407 401 410 0 nenh l=2e-06 w=8e-06 

m1033 414 416 415 0 nenh l=2e-06 w=8e-06 

m1034 415 418 417 0 nenh l=2e-06 w=6e-06 

m1035 417 271 419 0 nenh l=2e-06 w=5e-06 

m1036 419 421 420 0 nenh l=2e-06 w=5e-06 

m1037 420 278 415 0 nenh l=2e-06 w=6e-06 

m1038 415 283 422 0 nenh l=2e-06 w=8e-06 

m1039 422 424 423 0 nenh l=2e-06 w=1e-05 

m1040 0 419 425 0 nenh l=2e-06 w=6e-06 

m1041 3 329 419 3 penh l=2e-06 w=1.6e-05 

m1042 419 425 3 3 penh l=8e-06 w=4e-06 

m1043 3 419 425 3 penh l=2e-06 w=1.6e-05 

m1044 3 427 426 3 penh l=2e-06 w=1.6e-05 

m1045 3 329 427 3 penh l=2e-06 w=1.6e-05 

m1046 427 426 3 3 penh l=8e-06 w=4e-06 

m1047 426 427 0 0 nenh l=2e-06 w=6e-06 

m1048 0 329 423 0 nenh l=2e-06 w=4e-06 

m1049 423 288 414 0 nenh l=2e-06 w=1e-05 

m1050 414 283 428 0 nenh l=2e-06 w=8e-06 

m1051 428 278 417 0 nenh l=2e-06 w=7e-06 

m1052 417 421 427 0 nenh l=2e-06 w=6e-06 

m1053 427 271 420 0 nenh l=2e-06 w=6e-06 

m1054 420 418 428 0 nenh l=2e-06 w=7e-06 

m1055 428 416 422 0 nenh l=2e-06 w=8e-06 

m1056 429 431 430 0 nenh l=2e-06 w=8e-06 

m1057 430 433 432 0 nenh l=2e-06 w=6e-06 

m1058 432 305 434 0 nenh l=2e-06 w=5e-06 

m1059 434 436 435 0 nenh l=2e-06 w=5e-06 

m1060 435 301 430 0 nenh l=2e-06 w=6e-06 

m1061 430 297 437 0 nenh l=2e-06 w=8e-06 

m1062 437 439 438 0 nenh l=2e-06 w=1e-05 

m1063 0 434 440 0 nenh l=2e-06 w=6e-06 

m1064 3 329 434 3 penh l=2e-06 w=1.6e-05 

m1065 434 440 3 3 penh l=8e-06 w=4e-06 

m1066 3 434 440 3 penh l=2e-06 w=1.6e-05 

m1067 3 442 441 3 penh l=2e-06 w=1.6e-05 

m1068 3 329 442 3 penh l=2e-06 w=1.6e-05 

m1069 442 441 3 3 penh l=8e-06 w=4e-06 

m1070 441 442 0 0 nenh l=2e-06 w=6e-06 

m1071 0 329 438 0 nenh l=2e-06 w=4e-06 

m1072 438 293 429 0 nenh l=2e-06 w=1e-05 

m1073 429 297 443 0 nenh l=2e-06 w=8e-06 

m1074 443 301 432 0 nenh l=2e-06 w=7e-06 

m1075 432 436 442 0 nenh l=2e-06 w=6e-06 

m1076 442 305 435 0 nenh l=2e-06 w=6e-06 

m1077 435 433 443 0 nenh l=2e-06 w=7e-06 

m1078 443 431 437 0 nenh l=2e-06 w=8e-06 

m1079 444 366 445 0 nenh l=2e-06 w=6e-06 

m1080 445 447 446 0 nenh l=2e-06 w=6e-06 

m1081 0 444 448 0 nenh l=2e-06 w=6e-06 

m1082 3 329 444 3 penh l=2e-06 w=1e-05 

m1083 444 448 3 3 penh l=8e-06 w=4e-06 

m1084 3 444 448 3 penh l=2e-06 w=1.6e-05 

m1085 3 449 325 3 penh l=2e-06 w=1.6e-05 

m1086 3 329 449 3 penh l=2e-06 w=1e-05 

m1087 449 325 3 3 penh l=8e-06 w=4e-06 

m1088 325 449 0 0 nenh l=2e-06 w=6e-06 

m1089 0 329 446 0 nenh l=2e-06 w=1.2e-05 

m1090 446 451 450 0 nenh l=2e-06 w=6e-06 

m1091 450 366 449 0 nenh l=2e-06 w=6e-06 

m1092 449 367 446 0 nenh l=2e-06 w=6e-06 

m1093 452 385 453 0 nenh l=2e-06 w=6e-06 

m1094 453 455 454 0 nenh l=2e-06 w=6e-06 

m1095 0 452 456 0 nenh l=2e-06 w=6e-06 

m1096 3 329 452 3 penh l=2e-06 w=1e-05 

m1097 452 456 3 3 penh l=8e-06 w=4e-06 

m1098 3 452 456 3 penh l=2e-06 w=1.6e-05 

m1099 3 457 333 3 penh l=2e-06 w=1.6e-05 

m1100 3 329 457 3 penh l=2e-06 w=1e-05 

m1101 457 333 3 3 penh l=8e-06 w=4e-06 

m1102 333 457 0 0 nenh l=2e-06 w=6e-06 

m1103 0 329 454 0 nenh l=2e-06 w=1.2e-05 

m1104 454 459 458 0 nenh l=2e-06 w=6e-06 

m1105 458 385 457 0 nenh l=2e-06 w=6e-06 

m1106 457 386 454 0 nenh l=2e-06 w=6e-06 

m1107 460 404 461 0 nenh l=2e-06 w=6e-06 

m1108 461 463 462 0 nenh l=2e-06 w=6e-06 

m1109 0 460 464 0 nenh l=2e-06 w=6e-06 

m1110 3 329 460 3 penh l=2e-06 w=1e-05 

m1111 460 464 3 3 penh l=8e-06 w=4e-06 

m1112 3 460 464 3 penh l=2e-06 w=1.6e-05 

m1113 3 465 339 3 penh l=2e-06 w=1.6e-05 

m1114 3 329 465 3 penh l=2e-06 w=1e-05 

m1115 465 339 3 3 penh l=8e-06 w=4e-06 

m1116 339 465 0 0 nenh l=2e-06 w=6e-06 

m1117 0 329 462 0 nenh l=2e-06 w=1.2e-05 

m1118 462 467 466 0 nenh l=2e-06 w=6e-06 

m1119 466 404 465 0 nenh l=2e-06 w=6e-06 

m1120 465 405 462 0 nenh l=2e-06 w=6e-06 

m1121 468 426 469 0 nenh l=2e-06 w=4e-06 

m1122 469 425 470 0 nenh l=2e-06 w=4e-06 

m1123 0 469 471 0 nenh l=2e-06 w=6e-06 

m1124 3 329 469 3 penh l=2e-06 w=1.6e-05 

m1125 469 471 3 3 penh l=8e-06 w=4e-06 

m1126 3 469 471 3 penh l=2e-06 w=1.6e-05 

m1127 3 473 472 3 penh l=2e-06 w=1.6e-05 

m1128 3 329 473 3 penh l=2e-06 w=1.6e-05 

m1129 473 472 3 3 penh l=8e-06 w=4e-06 

m1130 472 473 0 0 nenh l=2e-06 w=6e-06 

m1131 0 329 474 0 nenh l=2e-06 w=4e-06 

m1132 474 441 468 0 nenh l=2e-06 w=8e-06 

m1133 468 425 473 0 nenh l=2e-06 w=4e-06 

m1134 473 426 470 0 nenh l=2e-06 w=4e-06 

m1135 470 440 474 0 nenh l=2e-06 w=8e-06 

m1136 475 456 476 0 nenh l=2e-06 w=8e-06 

m1137 476 471 477 0 nenh l=2e-06 w=6e-06 

m1138 477 325 478 0 nenh l=2e-06 w=5e-06 

m1139 478 448 479 0 nenh l=2e-06 w=5e-06 

m1140 479 472 476 0 nenh l=2e-06 w=6e-06 

m1141 476 333 480 0 nenh l=2e-06 w=8e-06 

m1142 480 464 481 0 nenh l=2e-06 w=1e-05 

m1143 0 478 351 0 nenh l=2e-06 w=6e-06 

m1144 3 329 478 3 penh l=2e-06 w=1.6e-05 

m1145 478 351 3 3 penh l=8e-06 w=4e-06 

m1146 3 478 351 3 penh l=2e-06 w=1.6e-05 

m1147 3 482 345 3 penh l=2e-06 w=1.6e-05 

m1148 3 329 482 3 penh l=2e-06 w=1.6e-05 

m1149 482 345 3 3 penh l=8e-06 w=4e-06 

m1150 345 482 0 0 nenh l=2e-06 w=6e-06 

m1151 0 329 481 0 nenh l=2e-06 w=4e-06 

m1152 481 339 475 0 nenh l=2e-06 w=1e-05 

m1153 475 333 483 0 nenh l=2e-06 w=8e-06 

m1154 483 472 477 0 nenh l=2e-06 w=7e-06 

m1155 477 448 482 0 nenh l=2e-06 w=6e-06 

m1156 482 325 479 0 nenh l=2e-06 w=6e-06 

m1157 479 471 483 0 nenh l=2e-06 w=7e-06 

m1158 483 456 480 0 nenh l=2e-06 w=8e-06 

m1159 484 486 485 0 nenh l=2e-06 w=1.2e-05 

m1160 484 488 487 0 nenh l=2e-06 w=1.2e-05 

m1161 487 490 489 0 nenh l=2e-06 w=1.2e-05 

m1162 489 492 491 0 nenh l=2e-06 w=1.4e-05 

m1163 0 485 447 0 nenh l=2e-06 w=6e-06 

m1164 3 329 485 3 penh l=2e-06 w=1e-05 

m1165 485 447 3 3 penh l=8e-06 w=4e-06 

m1166 3 485 447 3 penh l=2e-06 w=1.6e-05 

m1167 3 493 451 3 penh l=2e-06 w=1.6e-05 

m1168 3 329 493 3 penh l=2e-06 w=1e-05 

m1169 493 451 3 3 penh l=8e-06 w=4e-06 

m1170 451 493 0 0 nenh l=2e-06 w=6e-06 

m1171 0 329 491 0 nenh l=2e-06 w=1.4e-05 

m1172 494 495 491 0 nenh l=2e-06 w=8e-06 

m1173 491 488 496 0 nenh l=2e-06 w=1e-05 

m1174 496 498 497 0 nenh l=2e-06 w=1e-05 

m1175 497 499 491 0 nenh l=2e-06 w=8e-06 

m1176 491 500 493 0 nenh l=2e-06 w=6e-06 

m1177 493 492 494 0 nenh l=2e-06 w=6e-06 

m1178 494 490 497 0 nenh l=2e-06 w=8e-06 

m1179 501 503 502 0 nenh l=2e-06 w=1.2e-05 

m1180 501 505 504 0 nenh l=2e-06 w=1.2e-05 

m1181 504 507 506 0 nenh l=2e-06 w=1.2e-05 

m1182 506 509 508 0 nenh l=2e-06 w=1.4e-05 

m1183 0 502 455 0 nenh l=2e-06 w=6e-06 

m1184 3 329 502 3 penh l=2e-06 w=1e-05 

m1185 502 455 3 3 penh l=8e-06 w=4e-06 

m1186 3 502 455 3 penh l=2e-06 w=1.6e-05 

m1187 3 510 459 3 penh l=2e-06 w=1.6e-05 

m1188 3 329 510 3 penh l=2e-06 w=1e-05 

m1189 510 459 3 3 penh l=8e-06 w=4e-06 

m1190 459 510 0 0 nenh l=2e-06 w=6e-06 

m1191 0 329 508 0 nenh l=2e-06 w=1.4e-05 

m1192 511 512 508 0 nenh l=2e-06 w=8e-06 

m1193 508 505 513 0 nenh l=2e-06 w=1e-05 

m1194 513 515 514 0 nenh l=2e-06 w=1e-05 

m1195 514 516 508 0 nenh l=2e-06 w=8e-06 

m1196 508 517 510 0 nenh l=2e-06 w=6e-06 

m1197 510 509 511 0 nenh l=2e-06 w=6e-06 

m1198 511 507 514 0 nenh l=2e-06 w=8e-06 

m1199 518 520 519 0 nenh l=2e-06 w=1.2e-05 

m1200 518 522 521 0 nenh l=2e-06 w=1.2e-05 

m1201 521 524 523 0 nenh l=2e-06 w=1.2e-05 

m1202 523 526 525 0 nenh l=2e-06 w=1.4e-05 

m1203 0 519 463 0 nenh l=2e-06 w=6e-06 

m1204 3 329 519 3 penh l=2e-06 w=1e-05 

m1205 519 463 3 3 penh l=8e-06 w=4e-06 

m1206 3 519 463 3 penh l=2e-06 w=1.6e-05 

m1207 3 527 467 3 penh l=2e-06 w=1.6e-05 

m1208 3 329 527 3 penh l=2e-06 w=1e-05 

m1209 527 467 3 3 penh l=8e-06 w=4e-06 

m1210 467 527 0 0 nenh l=2e-06 w=6e-06 

m1211 0 329 525 0 nenh l=2e-06 w=1.4e-05 

m1212 528 529 525 0 nenh l=2e-06 w=8e-06 

m1213 525 522 530 0 nenh l=2e-06 w=1e-05 

m1214 530 532 531 0 nenh l=2e-06 w=1e-05 

m1215 531 533 525 0 nenh l=2e-06 w=8e-06 

m1216 525 534 527 0 nenh l=2e-06 w=6e-06 

m1217 527 526 528 0 nenh l=2e-06 w=6e-06 

m1218 528 524 531 0 nenh l=2e-06 w=8e-06 

m1219 535 327 536 3 penh l=2e-06 w=5e-06 

m1220 536 329 537 3 penh l=2e-06 w=5e-06 

m1221 537 538 3 3 penh l=2e-06 w=5e-06 

m1222 3 536 538 3 penh l=2e-06 w=6e-06 

m1223 538 28 3 3 penh l=2e-06 w=6e-06 

m1224 3 538 271 3 penh l=2e-06 w=2.5e-05 

m1225 535 329 536 0 nenh l=2e-06 w=5e-06 

m1226 536 327 539 0 nenh l=2e-06 w=5e-06 

m1227 539 538 0 0 nenh l=2e-06 w=5e-06 

m1228 0 536 540 0 nenh l=2e-06 w=1.3e-05 

m1229 540 28 538 0 nenh l=2e-06 w=1.2e-05 

m1230 0 538 271 0 nenh l=2e-06 w=1.4e-05 

m1231 541 223 542 0 nenh l=2e-06 w=8e-06 

m1232 542 544 543 0 nenh l=2e-06 w=6e-06 

m1233 543 228 541 0 nenh l=2e-06 w=8e-06 

m1234 541 546 545 0 nenh l=2e-06 w=1e-05 

m1235 0 542 403 0 nenh l=2e-06 w=6e-06 

m1236 403 542 3 3 penh l=2e-06 w=1.6e-05 

m1237 3 403 542 3 penh l=8e-06 w=4e-06 

m1238 542 329 3 3 penh l=2e-06 w=1e-05 

m1239 3 547 413 3 penh l=2e-06 w=1.6e-05 

m1240 3 413 547 3 penh l=8e-06 w=4e-06 

m1241 547 329 3 3 penh l=2e-06 w=1e-05 

m1242 413 547 0 0 nenh l=2e-06 w=6e-06 

m1243 0 329 545 0 nenh l=2e-06 w=1.4e-05 

m1244 545 549 548 0 nenh l=2e-06 w=1e-05 

m1245 548 228 542 0 nenh l=2e-06 w=8e-06 

m1246 542 551 550 0 nenh l=2e-06 w=6e-06 

m1247 550 223 548 0 nenh l=2e-06 w=8e-06 

m1248 543 551 547 0 nenh l=2e-06 w=6e-06 

m1249 547 544 550 0 nenh l=2e-06 w=6e-06 

m1250 552 549 553 0 nenh l=2e-06 w=8e-06 

m1251 553 223 554 0 nenh l=2e-06 w=4e-06 

m1252 554 546 552 0 nenh l=2e-06 w=8e-06 

m1253 552 551 555 0 nenh l=2e-06 w=1e-05 

m1254 0 553 421 0 nenh l=2e-06 w=6e-06 

m1255 3 329 553 3 penh l=2e-06 w=1e-05 

m1256 553 421 3 3 penh l=8e-06 w=4e-06 

m1257 3 553 421 3 penh l=2e-06 w=1.6e-05 

m1258 3 556 535 3 penh l=2e-06 w=1.6e-05 

m1259 3 329 556 3 penh l=2e-06 w=1e-05 

m1260 556 535 3 3 penh l=8e-06 w=4e-06 

m1261 535 556 0 0 nenh l=2e-06 w=6e-06 

m1262 0 329 555 0 nenh l=2e-06 w=1.4e-05 

m1263 555 544 557 0 nenh l=2e-06 w=1.2e-05 

m1264 557 549 554 0 nenh l=2e-06 w=6e-06 

m1265 554 228 556 0 nenh l=2e-06 w=4e-06 

m1266 556 546 557 0 nenh l=2e-06 w=6e-06 

m1267 558 551 559 0 nenh l=2e-06 w=8e-06 

m1268 559 546 560 0 nenh l=2e-06 w=6e-06 

m1269 560 544 558 0 nenh l=2e-06 w=8e-06 

m1270 558 228 561 0 nenh l=2e-06 w=1e-05 

m1271 0 559 384 0 nenh l=2e-06 w=6e-06 

m1272 3 329 559 3 penh l=2e-06 w=1e-05 

m1273 559 384 3 3 penh l=8e-06 w=4e-06 

m1274 3 559 384 3 penh l=2e-06 w=1.6e-05 

m1275 3 562 394 3 penh l=2e-06 w=1.6e-05 

m1276 3 329 562 3 penh l=2e-06 w=1e-05 

m1277 562 394 3 3 penh l=8e-06 w=4e-06 

m1278 394 562 0 0 nenh l=2e-06 w=6e-06 

m1279 0 329 561 0 nenh l=2e-06 w=1.4e-05 

m1280 561 223 563 0 nenh l=2e-06 w=1e-05 

m1281 563 544 559 0 nenh l=2e-06 w=8e-06 

m1282 559 549 564 0 nenh l=2e-06 w=6e-06 

m1283 564 551 563 0 nenh l=2e-06 w=8e-06 

m1284 560 549 562 0 nenh l=2e-06 w=6e-06 

m1285 562 546 564 0 nenh l=2e-06 w=6e-06 

m1286 565 549 566 0 nenh l=2e-06 w=8e-06 

m1287 566 228 567 0 nenh l=2e-06 w=6e-06 

m1288 567 546 565 0 nenh l=2e-06 w=8e-06 

m1289 565 544 568 0 nenh l=2e-06 w=1e-05 

m1290 0 566 365 0 nenh l=2e-06 w=6e-06 

m1291 365 566 3 3 penh l=2e-06 w=1.6e-05 

m1292 3 365 566 3 penh l=8e-06 w=4e-06 

m1293 566 329 3 3 penh l=2e-06 w=1e-05 

m1294 3 569 375 3 penh l=2e-06 w=1.6e-05 

m1295 3 375 569 3 penh l=8e-06 w=4e-06 

m1296 569 329 3 3 penh l=2e-06 w=1e-05 

m1297 375 569 0 0 nenh l=2e-06 w=6e-06 

m1298 0 329 568 0 nenh l=2e-06 w=1.4e-05 

m1299 568 551 570 0 nenh l=2e-06 w=1e-05 

m1300 570 546 566 0 nenh l=2e-06 w=8e-06 

m1301 566 223 571 0 nenh l=2e-06 w=6e-06 

m1302 571 549 570 0 nenh l=2e-06 w=8e-06 

m1303 567 223 569 0 nenh l=2e-06 w=6e-06 

m1304 569 228 571 0 nenh l=2e-06 w=6e-06 

m1305 572 327 573 3 penh l=2e-06 w=5e-06 

m1306 573 329 574 3 penh l=2e-06 w=5e-06 

m1307 574 575 3 3 penh l=2e-06 w=5e-06 

m1308 3 573 575 3 penh l=2e-06 w=6e-06 

m1309 575 28 3 3 penh l=2e-06 w=6e-06 

m1310 3 575 278 3 penh l=2e-06 w=2.5e-05 

m1311 572 329 573 0 nenh l=2e-06 w=5e-06 

m1312 573 327 576 0 nenh l=2e-06 w=5e-06 

m1313 576 575 0 0 nenh l=2e-06 w=5e-06 

m1314 0 573 577 0 nenh l=2e-06 w=1.3e-05 

m1315 577 28 575 0 nenh l=2e-06 w=1.2e-05 

m1316 0 575 278 0 nenh l=2e-06 w=1.4e-05 

m1317 578 204 579 0 nenh l=2e-06 w=8e-06 

m1318 579 581 580 0 nenh l=2e-06 w=6e-06 

m1319 580 209 578 0 nenh l=2e-06 w=8e-06 

m1320 578 583 582 0 nenh l=2e-06 w=1e-05 

m1321 0 579 401 0 nenh l=2e-06 w=6e-06 

m1322 401 579 3 3 penh l=2e-06 w=1.6e-05 

m1323 3 401 579 3 penh l=8e-06 w=4e-06 

m1324 579 329 3 3 penh l=2e-06 w=1e-05 

m1325 3 584 408 3 penh l=2e-06 w=1.6e-05 

m1326 3 408 584 3 penh l=8e-06 w=4e-06 

m1327 584 329 3 3 penh l=2e-06 w=1e-05 

m1328 408 584 0 0 nenh l=2e-06 w=6e-06 

m1329 0 329 582 0 nenh l=2e-06 w=1.4e-05 

m1330 582 586 585 0 nenh l=2e-06 w=1e-05 

m1331 585 209 579 0 nenh l=2e-06 w=8e-06 

m1332 579 588 587 0 nenh l=2e-06 w=6e-06 

m1333 587 204 585 0 nenh l=2e-06 w=8e-06 

m1334 580 588 584 0 nenh l=2e-06 w=6e-06 

m1335 584 581 587 0 nenh l=2e-06 w=6e-06 

m1336 589 586 590 0 nenh l=2e-06 w=8e-06 

m1337 590 204 591 0 nenh l=2e-06 w=4e-06 

m1338 591 583 589 0 nenh l=2e-06 w=8e-06 

m1339 589 588 592 0 nenh l=2e-06 w=1e-05 

m1340 0 590 418 0 nenh l=2e-06 w=6e-06 

m1341 3 329 590 3 penh l=2e-06 w=1e-05 

m1342 590 418 3 3 penh l=8e-06 w=4e-06 

m1343 3 590 418 3 penh l=2e-06 w=1.6e-05 

m1344 3 593 572 3 penh l=2e-06 w=1.6e-05 

m1345 3 329 593 3 penh l=2e-06 w=1e-05 

m1346 593 572 3 3 penh l=8e-06 w=4e-06 

m1347 572 593 0 0 nenh l=2e-06 w=6e-06 

m1348 0 329 592 0 nenh l=2e-06 w=1.4e-05 

m1349 592 581 594 0 nenh l=2e-06 w=1.2e-05 

m1350 594 586 591 0 nenh l=2e-06 w=6e-06 

m1351 591 209 593 0 nenh l=2e-06 w=4e-06 

m1352 593 583 594 0 nenh l=2e-06 w=6e-06 

m1353 595 588 596 0 nenh l=2e-06 w=8e-06 

m1354 596 583 597 0 nenh l=2e-06 w=6e-06 

m1355 597 581 595 0 nenh l=2e-06 w=8e-06 

m1356 595 209 598 0 nenh l=2e-06 w=1e-05 

m1357 0 596 382 0 nenh l=2e-06 w=6e-06 

m1358 3 329 596 3 penh l=2e-06 w=1e-05 

m1359 596 382 3 3 penh l=8e-06 w=4e-06 

m1360 3 596 382 3 penh l=2e-06 w=1.6e-05 

m1361 3 599 389 3 penh l=2e-06 w=1.6e-05 

m1362 3 329 599 3 penh l=2e-06 w=1e-05 

m1363 599 389 3 3 penh l=8e-06 w=4e-06 

m1364 389 599 0 0 nenh l=2e-06 w=6e-06 

m1365 0 329 598 0 nenh l=2e-06 w=1.4e-05 

m1366 598 204 600 0 nenh l=2e-06 w=1e-05 

m1367 600 581 596 0 nenh l=2e-06 w=8e-06 

m1368 596 586 601 0 nenh l=2e-06 w=6e-06 

m1369 601 588 600 0 nenh l=2e-06 w=8e-06 

m1370 597 586 599 0 nenh l=2e-06 w=6e-06 

m1371 599 583 601 0 nenh l=2e-06 w=6e-06 

m1372 602 586 603 0 nenh l=2e-06 w=8e-06 

m1373 603 209 604 0 nenh l=2e-06 w=6e-06 

m1374 604 583 602 0 nenh l=2e-06 w=8e-06 

m1375 602 581 605 0 nenh l=2e-06 w=1e-05 

m1376 0 603 363 0 nenh l=2e-06 w=6e-06 

m1377 363 603 3 3 penh l=2e-06 w=1.6e-05 

m1378 3 363 603 3 penh l=8e-06 w=4e-06 

m1379 603 329 3 3 penh l=2e-06 w=1e-05 

m1380 3 606 370 3 penh l=2e-06 w=1.6e-05 

m1381 3 370 606 3 penh l=8e-06 w=4e-06 

m1382 606 329 3 3 penh l=2e-06 w=1e-05 

m1383 370 606 0 0 nenh l=2e-06 w=6e-06 

m1384 0 329 605 0 nenh l=2e-06 w=1.4e-05 

m1385 605 588 607 0 nenh l=2e-06 w=1e-05 

m1386 607 583 603 0 nenh l=2e-06 w=8e-06 

m1387 603 204 608 0 nenh l=2e-06 w=6e-06 

m1388 608 586 607 0 nenh l=2e-06 w=8e-06 

m1389 604 204 606 0 nenh l=2e-06 w=6e-06 

m1390 606 209 608 0 nenh l=2e-06 w=6e-06 

m1391 609 327 610 3 penh l=2e-06 w=5e-06 

m1392 610 329 611 3 penh l=2e-06 w=5e-06 

m1393 611 612 3 3 penh l=2e-06 w=5e-06 

m1394 3 610 612 3 penh l=2e-06 w=6e-06 

m1395 612 28 3 3 penh l=2e-06 w=6e-06 

m1396 3 612 283 3 penh l=2e-06 w=2.5e-05 

m1397 609 329 610 0 nenh l=2e-06 w=5e-06 

m1398 610 327 613 0 nenh l=2e-06 w=5e-06 

m1399 613 612 0 0 nenh l=2e-06 w=5e-06 

m1400 0 610 614 0 nenh l=2e-06 w=1.3e-05 

m1401 614 28 612 0 nenh l=2e-06 w=1.2e-05 

m1402 0 612 283 0 nenh l=2e-06 w=1.4e-05 

m1403 615 185 616 0 nenh l=2e-06 w=8e-06 

m1404 616 618 617 0 nenh l=2e-06 w=6e-06 

m1405 617 190 615 0 nenh l=2e-06 w=8e-06 

m1406 615 620 619 0 nenh l=2e-06 w=1e-05 

m1407 0 616 399 0 nenh l=2e-06 w=6e-06 

m1408 399 616 3 3 penh l=2e-06 w=1.6e-05 

m1409 3 399 616 3 penh l=8e-06 w=4e-06 

m1410 616 329 3 3 penh l=2e-06 w=1e-05 

m1411 3 621 412 3 penh l=2e-06 w=1.6e-05 

m1412 3 412 621 3 penh l=8e-06 w=4e-06 

m1413 621 329 3 3 penh l=2e-06 w=1e-05 

m1414 412 621 0 0 nenh l=2e-06 w=6e-06 

m1415 0 329 619 0 nenh l=2e-06 w=1.4e-05 

m1416 619 623 622 0 nenh l=2e-06 w=1e-05 

m1417 622 190 616 0 nenh l=2e-06 w=8e-06 

m1418 616 625 624 0 nenh l=2e-06 w=6e-06 

m1419 624 185 622 0 nenh l=2e-06 w=8e-06 

m1420 617 625 621 0 nenh l=2e-06 w=6e-06 

m1421 621 618 624 0 nenh l=2e-06 w=6e-06 

m1422 626 623 627 0 nenh l=2e-06 w=8e-06 

m1423 627 185 628 0 nenh l=2e-06 w=4e-06 

m1424 628 620 626 0 nenh l=2e-06 w=8e-06 

m1425 626 625 629 0 nenh l=2e-06 w=1e-05 

m1426 0 627 416 0 nenh l=2e-06 w=6e-06 

m1427 3 329 627 3 penh l=2e-06 w=1e-05 

m1428 627 416 3 3 penh l=8e-06 w=4e-06 

m1429 3 627 416 3 penh l=2e-06 w=1.6e-05 

m1430 3 630 609 3 penh l=2e-06 w=1.6e-05 

m1431 3 329 630 3 penh l=2e-06 w=1e-05 

m1432 630 609 3 3 penh l=8e-06 w=4e-06 

m1433 609 630 0 0 nenh l=2e-06 w=6e-06 

m1434 0 329 629 0 nenh l=2e-06 w=1.4e-05 

m1435 629 618 631 0 nenh l=2e-06 w=1.2e-05 

m1436 631 623 628 0 nenh l=2e-06 w=6e-06 

m1437 628 190 630 0 nenh l=2e-06 w=4e-06 

m1438 630 620 631 0 nenh l=2e-06 w=6e-06 

m1439 632 625 633 0 nenh l=2e-06 w=8e-06 

m1440 633 620 634 0 nenh l=2e-06 w=6e-06 

m1441 634 618 632 0 nenh l=2e-06 w=8e-06 

m1442 632 190 635 0 nenh l=2e-06 w=1e-05 

m1443 0 633 380 0 nenh l=2e-06 w=6e-06 

m1444 3 329 633 3 penh l=2e-06 w=1e-05 

m1445 633 380 3 3 penh l=8e-06 w=4e-06 

m1446 3 633 380 3 penh l=2e-06 w=1.6e-05 

m1447 3 636 393 3 penh l=2e-06 w=1.6e-05 

m1448 3 329 636 3 penh l=2e-06 w=1e-05 

m1449 636 393 3 3 penh l=8e-06 w=4e-06 

m1450 393 636 0 0 nenh l=2e-06 w=6e-06 

m1451 0 329 635 0 nenh l=2e-06 w=1.4e-05 

m1452 635 185 637 0 nenh l=2e-06 w=1e-05 

m1453 637 618 633 0 nenh l=2e-06 w=8e-06 

m1454 633 623 638 0 nenh l=2e-06 w=6e-06 

m1455 638 625 637 0 nenh l=2e-06 w=8e-06 

m1456 634 623 636 0 nenh l=2e-06 w=6e-06 

m1457 636 620 638 0 nenh l=2e-06 w=6e-06 

m1458 639 623 640 0 nenh l=2e-06 w=8e-06 

m1459 640 190 641 0 nenh l=2e-06 w=6e-06 

m1460 641 620 639 0 nenh l=2e-06 w=8e-06 

m1461 639 618 642 0 nenh l=2e-06 w=1e-05 

m1462 0 640 361 0 nenh l=2e-06 w=6e-06 

m1463 361 640 3 3 penh l=2e-06 w=1.6e-05 

m1464 3 361 640 3 penh l=8e-06 w=4e-06 

m1465 640 329 3 3 penh l=2e-06 w=1e-05 

m1466 3 643 374 3 penh l=2e-06 w=1.6e-05 

m1467 3 374 643 3 penh l=8e-06 w=4e-06 

m1468 643 329 3 3 penh l=2e-06 w=1e-05 

m1469 374 643 0 0 nenh l=2e-06 w=6e-06 

m1470 0 329 642 0 nenh l=2e-06 w=1.4e-05 

m1471 642 625 644 0 nenh l=2e-06 w=1e-05 

m1472 644 620 640 0 nenh l=2e-06 w=8e-06 

m1473 640 185 645 0 nenh l=2e-06 w=6e-06 

m1474 645 623 644 0 nenh l=2e-06 w=8e-06 

m1475 641 185 643 0 nenh l=2e-06 w=6e-06 

m1476 643 190 645 0 nenh l=2e-06 w=6e-06 

m1477 646 327 647 3 penh l=2e-06 w=5e-06 

m1478 647 329 648 3 penh l=2e-06 w=5e-06 

m1479 648 649 3 3 penh l=2e-06 w=5e-06 

m1480 3 647 649 3 penh l=2e-06 w=6e-06 

m1481 649 28 3 3 penh l=2e-06 w=6e-06 

m1482 3 649 288 3 penh l=2e-06 w=2.5e-05 

m1483 646 329 647 0 nenh l=2e-06 w=5e-06 

m1484 647 327 650 0 nenh l=2e-06 w=5e-06 

m1485 650 649 0 0 nenh l=2e-06 w=5e-06 

m1486 0 647 651 0 nenh l=2e-06 w=1.3e-05 

m1487 651 28 649 0 nenh l=2e-06 w=1.2e-05 

m1488 0 649 288 0 nenh l=2e-06 w=1.4e-05 

m1489 652 166 653 0 nenh l=2e-06 w=8e-06 

m1490 653 655 654 0 nenh l=2e-06 w=6e-06 

m1491 654 171 652 0 nenh l=2e-06 w=8e-06 

m1492 652 657 656 0 nenh l=2e-06 w=1e-05 

m1493 0 653 397 0 nenh l=2e-06 w=6e-06 

m1494 397 653 3 3 penh l=2e-06 w=1.6e-05 

m1495 3 397 653 3 penh l=8e-06 w=4e-06 

m1496 653 329 3 3 penh l=2e-06 w=1e-05 

m1497 3 658 411 3 penh l=2e-06 w=1.6e-05 

m1498 3 411 658 3 penh l=8e-06 w=4e-06 

m1499 658 329 3 3 penh l=2e-06 w=1e-05 

m1500 411 658 0 0 nenh l=2e-06 w=6e-06 

m1501 0 329 656 0 nenh l=2e-06 w=1.4e-05 

m1502 656 660 659 0 nenh l=2e-06 w=1e-05 

m1503 659 171 653 0 nenh l=2e-06 w=8e-06 

m1504 653 662 661 0 nenh l=2e-06 w=6e-06 

m1505 661 166 659 0 nenh l=2e-06 w=8e-06 

m1506 654 662 658 0 nenh l=2e-06 w=6e-06 

m1507 658 655 661 0 nenh l=2e-06 w=6e-06 

m1508 663 660 664 0 nenh l=2e-06 w=8e-06 

m1509 664 166 665 0 nenh l=2e-06 w=4e-06 

m1510 665 657 663 0 nenh l=2e-06 w=8e-06 

m1511 663 662 666 0 nenh l=2e-06 w=1e-05 

m1512 0 664 424 0 nenh l=2e-06 w=6e-06 

m1513 3 329 664 3 penh l=2e-06 w=1e-05 

m1514 664 424 3 3 penh l=8e-06 w=4e-06 

m1515 3 664 424 3 penh l=2e-06 w=1.6e-05 

m1516 3 667 646 3 penh l=2e-06 w=1.6e-05 

m1517 3 329 667 3 penh l=2e-06 w=1e-05 

m1518 667 646 3 3 penh l=8e-06 w=4e-06 

m1519 646 667 0 0 nenh l=2e-06 w=6e-06 

m1520 0 329 666 0 nenh l=2e-06 w=1.4e-05 

m1521 666 655 668 0 nenh l=2e-06 w=1.2e-05 

m1522 668 660 665 0 nenh l=2e-06 w=6e-06 

m1523 665 171 667 0 nenh l=2e-06 w=4e-06 

m1524 667 657 668 0 nenh l=2e-06 w=6e-06 

m1525 669 662 670 0 nenh l=2e-06 w=8e-06 

m1526 670 657 671 0 nenh l=2e-06 w=6e-06 

m1527 671 655 669 0 nenh l=2e-06 w=8e-06 

m1528 669 171 672 0 nenh l=2e-06 w=1e-05 

m1529 0 670 378 0 nenh l=2e-06 w=6e-06 

m1530 3 329 670 3 penh l=2e-06 w=1e-05 

m1531 670 378 3 3 penh l=8e-06 w=4e-06 

m1532 3 670 378 3 penh l=2e-06 w=1.6e-05 

m1533 3 673 392 3 penh l=2e-06 w=1.6e-05 

m1534 3 329 673 3 penh l=2e-06 w=1e-05 

m1535 673 392 3 3 penh l=8e-06 w=4e-06 

m1536 392 673 0 0 nenh l=2e-06 w=6e-06 

m1537 0 329 672 0 nenh l=2e-06 w=1.4e-05 

m1538 672 166 674 0 nenh l=2e-06 w=1e-05 

m1539 674 655 670 0 nenh l=2e-06 w=8e-06 

m1540 670 660 675 0 nenh l=2e-06 w=6e-06 

m1541 675 662 674 0 nenh l=2e-06 w=8e-06 

m1542 671 660 673 0 nenh l=2e-06 w=6e-06 

m1543 673 657 675 0 nenh l=2e-06 w=6e-06 

m1544 676 660 677 0 nenh l=2e-06 w=8e-06 

m1545 677 171 678 0 nenh l=2e-06 w=6e-06 

m1546 678 657 676 0 nenh l=2e-06 w=8e-06 

m1547 676 655 679 0 nenh l=2e-06 w=1e-05 

m1548 0 677 359 0 nenh l=2e-06 w=6e-06 

m1549 359 677 3 3 penh l=2e-06 w=1.6e-05 

m1550 3 359 677 3 penh l=8e-06 w=4e-06 

m1551 677 329 3 3 penh l=2e-06 w=1e-05 

m1552 3 680 373 3 penh l=2e-06 w=1.6e-05 

m1553 3 373 680 3 penh l=8e-06 w=4e-06 

m1554 680 329 3 3 penh l=2e-06 w=1e-05 

m1555 373 680 0 0 nenh l=2e-06 w=6e-06 

m1556 0 329 679 0 nenh l=2e-06 w=1.4e-05 

m1557 679 662 681 0 nenh l=2e-06 w=1e-05 

m1558 681 657 677 0 nenh l=2e-06 w=8e-06 

m1559 677 166 682 0 nenh l=2e-06 w=6e-06 

m1560 682 660 681 0 nenh l=2e-06 w=8e-06 

m1561 678 166 680 0 nenh l=2e-06 w=6e-06 

m1562 680 171 682 0 nenh l=2e-06 w=6e-06 

m1563 683 327 684 3 penh l=2e-06 w=5e-06 

m1564 684 329 685 3 penh l=2e-06 w=5e-06 

m1565 685 686 3 3 penh l=2e-06 w=5e-06 

m1566 3 684 686 3 penh l=2e-06 w=6e-06 

m1567 686 28 3 3 penh l=2e-06 w=6e-06 

m1568 3 686 293 3 penh l=2e-06 w=2.5e-05 

m1569 683 329 684 0 nenh l=2e-06 w=5e-06 

m1570 684 327 687 0 nenh l=2e-06 w=5e-06 

m1571 687 686 0 0 nenh l=2e-06 w=5e-06 

m1572 0 684 688 0 nenh l=2e-06 w=1.3e-05 

m1573 688 28 686 0 nenh l=2e-06 w=1.2e-05 

m1574 0 686 293 0 nenh l=2e-06 w=1.4e-05 

m1575 689 146 690 0 nenh l=2e-06 w=8e-06 

m1576 690 692 691 0 nenh l=2e-06 w=6e-06 

m1577 691 151 689 0 nenh l=2e-06 w=8e-06 

m1578 689 694 693 0 nenh l=2e-06 w=1e-05 

m1579 0 690 520 0 nenh l=2e-06 w=6e-06 

m1580 520 690 3 3 penh l=2e-06 w=1.6e-05 

m1581 3 520 690 3 penh l=8e-06 w=4e-06 

m1582 690 329 3 3 penh l=2e-06 w=1e-05 

m1583 3 695 532 3 penh l=2e-06 w=1.6e-05 

m1584 3 532 695 3 penh l=8e-06 w=4e-06 

m1585 695 329 3 3 penh l=2e-06 w=1e-05 

m1586 532 695 0 0 nenh l=2e-06 w=6e-06 

m1587 0 329 693 0 nenh l=2e-06 w=1.4e-05 

m1588 693 697 696 0 nenh l=2e-06 w=1e-05 

m1589 696 151 690 0 nenh l=2e-06 w=8e-06 

m1590 690 699 698 0 nenh l=2e-06 w=6e-06 

m1591 698 146 696 0 nenh l=2e-06 w=8e-06 

m1592 691 699 695 0 nenh l=2e-06 w=6e-06 

m1593 695 692 698 0 nenh l=2e-06 w=6e-06 

m1594 700 697 701 0 nenh l=2e-06 w=8e-06 

m1595 701 146 702 0 nenh l=2e-06 w=4e-06 

m1596 702 694 700 0 nenh l=2e-06 w=8e-06 

m1597 700 699 703 0 nenh l=2e-06 w=1e-05 

m1598 0 701 439 0 nenh l=2e-06 w=6e-06 

m1599 3 329 701 3 penh l=2e-06 w=1e-05 

m1600 701 439 3 3 penh l=8e-06 w=4e-06 

m1601 3 701 439 3 penh l=2e-06 w=1.6e-05 

m1602 3 704 683 3 penh l=2e-06 w=1.6e-05 

m1603 3 329 704 3 penh l=2e-06 w=1e-05 

m1604 704 683 3 3 penh l=8e-06 w=4e-06 

m1605 683 704 0 0 nenh l=2e-06 w=6e-06 

m1606 0 329 703 0 nenh l=2e-06 w=1.4e-05 

m1607 703 692 705 0 nenh l=2e-06 w=1.2e-05 

m1608 705 697 702 0 nenh l=2e-06 w=6e-06 

m1609 702 151 704 0 nenh l=2e-06 w=4e-06 

m1610 704 694 705 0 nenh l=2e-06 w=6e-06 

m1611 706 699 707 0 nenh l=2e-06 w=8e-06 

m1612 707 694 708 0 nenh l=2e-06 w=6e-06 

m1613 708 692 706 0 nenh l=2e-06 w=8e-06 

m1614 706 151 709 0 nenh l=2e-06 w=1e-05 

m1615 0 707 503 0 nenh l=2e-06 w=6e-06 

m1616 3 329 707 3 penh l=2e-06 w=1e-05 

m1617 707 503 3 3 penh l=8e-06 w=4e-06 

m1618 3 707 503 3 penh l=2e-06 w=1.6e-05 

m1619 3 710 515 3 penh l=2e-06 w=1.6e-05 

m1620 3 329 710 3 penh l=2e-06 w=1e-05 

m1621 710 515 3 3 penh l=8e-06 w=4e-06 

m1622 515 710 0 0 nenh l=2e-06 w=6e-06 

m1623 0 329 709 0 nenh l=2e-06 w=1.4e-05 

m1624 709 146 711 0 nenh l=2e-06 w=1e-05 

m1625 711 692 707 0 nenh l=2e-06 w=8e-06 

m1626 707 697 712 0 nenh l=2e-06 w=6e-06 

m1627 712 699 711 0 nenh l=2e-06 w=8e-06 

m1628 708 697 710 0 nenh l=2e-06 w=6e-06 

m1629 710 694 712 0 nenh l=2e-06 w=6e-06 

m1630 713 697 714 0 nenh l=2e-06 w=8e-06 

m1631 714 151 715 0 nenh l=2e-06 w=6e-06 

m1632 715 694 713 0 nenh l=2e-06 w=8e-06 

m1633 713 692 716 0 nenh l=2e-06 w=1e-05 

m1634 0 714 490 0 nenh l=2e-06 w=6e-06 

m1635 490 714 3 3 penh l=2e-06 w=1.6e-05 

m1636 3 490 714 3 penh l=8e-06 w=4e-06 

m1637 714 329 3 3 penh l=2e-06 w=1e-05 

m1638 3 717 495 3 penh l=2e-06 w=1.6e-05 

m1639 3 495 717 3 penh l=8e-06 w=4e-06 

m1640 717 329 3 3 penh l=2e-06 w=1e-05 

m1641 495 717 0 0 nenh l=2e-06 w=6e-06 

m1642 0 329 716 0 nenh l=2e-06 w=1.4e-05 

m1643 716 699 718 0 nenh l=2e-06 w=1e-05 

m1644 718 694 714 0 nenh l=2e-06 w=8e-06 

m1645 714 146 719 0 nenh l=2e-06 w=6e-06 

m1646 719 697 718 0 nenh l=2e-06 w=8e-06 

m1647 715 146 717 0 nenh l=2e-06 w=6e-06 

m1648 717 151 719 0 nenh l=2e-06 w=6e-06 

m1649 720 327 721 3 penh l=2e-06 w=5e-06 

m1650 721 329 722 3 penh l=2e-06 w=5e-06 

m1651 722 723 3 3 penh l=2e-06 w=5e-06 

m1652 3 721 723 3 penh l=2e-06 w=6e-06 

m1653 723 28 3 3 penh l=2e-06 w=6e-06 

m1654 3 723 297 3 penh l=2e-06 w=2.5e-05 

m1655 720 329 721 0 nenh l=2e-06 w=5e-06 

m1656 721 327 724 0 nenh l=2e-06 w=5e-06 

m1657 724 723 0 0 nenh l=2e-06 w=5e-06 

m1658 0 721 725 0 nenh l=2e-06 w=1.3e-05 

m1659 725 28 723 0 nenh l=2e-06 w=1.2e-05 

m1660 0 723 297 0 nenh l=2e-06 w=1.4e-05 

m1661 726 126 727 0 nenh l=2e-06 w=8e-06 

m1662 727 729 728 0 nenh l=2e-06 w=6e-06 

m1663 728 131 726 0 nenh l=2e-06 w=8e-06 

m1664 726 731 730 0 nenh l=2e-06 w=1e-05 

m1665 0 727 522 0 nenh l=2e-06 w=6e-06 

m1666 522 727 3 3 penh l=2e-06 w=1.6e-05 

m1667 3 522 727 3 penh l=8e-06 w=4e-06 

m1668 727 329 3 3 penh l=2e-06 w=1e-05 

m1669 3 732 533 3 penh l=2e-06 w=1.6e-05 

m1670 3 533 732 3 penh l=8e-06 w=4e-06 

m1671 732 329 3 3 penh l=2e-06 w=1e-05 

m1672 533 732 0 0 nenh l=2e-06 w=6e-06 

m1673 0 329 730 0 nenh l=2e-06 w=1.4e-05 

m1674 730 734 733 0 nenh l=2e-06 w=1e-05 

m1675 733 131 727 0 nenh l=2e-06 w=8e-06 

m1676 727 736 735 0 nenh l=2e-06 w=6e-06 

m1677 735 126 733 0 nenh l=2e-06 w=8e-06 

m1678 728 736 732 0 nenh l=2e-06 w=6e-06 

m1679 732 729 735 0 nenh l=2e-06 w=6e-06 

m1680 737 734 738 0 nenh l=2e-06 w=8e-06 

m1681 738 126 739 0 nenh l=2e-06 w=4e-06 

m1682 739 731 737 0 nenh l=2e-06 w=8e-06 

m1683 737 736 740 0 nenh l=2e-06 w=1e-05 

m1684 0 738 431 0 nenh l=2e-06 w=6e-06 

m1685 3 329 738 3 penh l=2e-06 w=1e-05 

m1686 738 431 3 3 penh l=8e-06 w=4e-06 

m1687 3 738 431 3 penh l=2e-06 w=1.6e-05 

m1688 3 741 720 3 penh l=2e-06 w=1.6e-05 

m1689 3 329 741 3 penh l=2e-06 w=1e-05 

m1690 741 720 3 3 penh l=8e-06 w=4e-06 

m1691 720 741 0 0 nenh l=2e-06 w=6e-06 

m1692 0 329 740 0 nenh l=2e-06 w=1.4e-05 

m1693 740 729 742 0 nenh l=2e-06 w=1.2e-05 

m1694 742 734 739 0 nenh l=2e-06 w=6e-06 

m1695 739 131 741 0 nenh l=2e-06 w=4e-06 

m1696 741 731 742 0 nenh l=2e-06 w=6e-06 

m1697 743 736 744 0 nenh l=2e-06 w=8e-06 

m1698 744 731 745 0 nenh l=2e-06 w=6e-06 

m1699 745 729 743 0 nenh l=2e-06 w=8e-06 

m1700 743 131 746 0 nenh l=2e-06 w=1e-05 

m1701 0 744 505 0 nenh l=2e-06 w=6e-06 

m1702 3 329 744 3 penh l=2e-06 w=1e-05 

m1703 744 505 3 3 penh l=8e-06 w=4e-06 

m1704 3 744 505 3 penh l=2e-06 w=1.6e-05 

m1705 3 747 516 3 penh l=2e-06 w=1.6e-05 

m1706 3 329 747 3 penh l=2e-06 w=1e-05 

m1707 747 516 3 3 penh l=8e-06 w=4e-06 

m1708 516 747 0 0 nenh l=2e-06 w=6e-06 

m1709 0 329 746 0 nenh l=2e-06 w=1.4e-05 

m1710 746 126 748 0 nenh l=2e-06 w=1e-05 

m1711 748 729 744 0 nenh l=2e-06 w=8e-06 

m1712 744 734 749 0 nenh l=2e-06 w=6e-06 

m1713 749 736 748 0 nenh l=2e-06 w=8e-06 

m1714 745 734 747 0 nenh l=2e-06 w=6e-06 

m1715 747 731 749 0 nenh l=2e-06 w=6e-06 

m1716 750 734 751 0 nenh l=2e-06 w=8e-06 

m1717 751 131 752 0 nenh l=2e-06 w=6e-06 

m1718 752 731 750 0 nenh l=2e-06 w=8e-06 

m1719 750 729 753 0 nenh l=2e-06 w=1e-05 

m1720 0 751 492 0 nenh l=2e-06 w=6e-06 

m1721 492 751 3 3 penh l=2e-06 w=1.6e-05 

m1722 3 492 751 3 penh l=8e-06 w=4e-06 

m1723 751 329 3 3 penh l=2e-06 w=1e-05 

m1724 3 754 500 3 penh l=2e-06 w=1.6e-05 

m1725 3 500 754 3 penh l=8e-06 w=4e-06 

m1726 754 329 3 3 penh l=2e-06 w=1e-05 

m1727 500 754 0 0 nenh l=2e-06 w=6e-06 

m1728 0 329 753 0 nenh l=2e-06 w=1.4e-05 

m1729 753 736 755 0 nenh l=2e-06 w=1e-05 

m1730 755 731 751 0 nenh l=2e-06 w=8e-06 

m1731 751 126 756 0 nenh l=2e-06 w=6e-06 

m1732 756 734 755 0 nenh l=2e-06 w=8e-06 

m1733 752 126 754 0 nenh l=2e-06 w=6e-06 

m1734 754 131 756 0 nenh l=2e-06 w=6e-06 

m1735 757 327 758 3 penh l=2e-06 w=5e-06 

m1736 758 329 759 3 penh l=2e-06 w=5e-06 

m1737 759 760 3 3 penh l=2e-06 w=5e-06 

m1738 3 758 760 3 penh l=2e-06 w=6e-06 

m1739 760 28 3 3 penh l=2e-06 w=6e-06 

m1740 3 760 301 3 penh l=2e-06 w=2.5e-05 

m1741 757 329 758 0 nenh l=2e-06 w=5e-06 

m1742 758 327 761 0 nenh l=2e-06 w=5e-06 

m1743 761 760 0 0 nenh l=2e-06 w=5e-06 

m1744 0 758 762 0 nenh l=2e-06 w=1.3e-05 

m1745 762 28 760 0 nenh l=2e-06 w=1.2e-05 

m1746 0 760 301 0 nenh l=2e-06 w=1.4e-05 

m1747 763 106 764 0 nenh l=2e-06 w=8e-06 

m1748 764 766 765 0 nenh l=2e-06 w=6e-06 

m1749 765 111 763 0 nenh l=2e-06 w=8e-06 

m1750 763 768 767 0 nenh l=2e-06 w=1e-05 

m1751 0 764 524 0 nenh l=2e-06 w=6e-06 

m1752 524 764 3 3 penh l=2e-06 w=1.6e-05 

m1753 3 524 764 3 penh l=8e-06 w=4e-06 

m1754 764 329 3 3 penh l=2e-06 w=1e-05 

m1755 3 769 529 3 penh l=2e-06 w=1.6e-05 

m1756 3 529 769 3 penh l=8e-06 w=4e-06 

m1757 769 329 3 3 penh l=2e-06 w=1e-05 

m1758 529 769 0 0 nenh l=2e-06 w=6e-06 

m1759 0 329 767 0 nenh l=2e-06 w=1.4e-05 

m1760 767 771 770 0 nenh l=2e-06 w=1e-05 

m1761 770 111 764 0 nenh l=2e-06 w=8e-06 

m1762 764 773 772 0 nenh l=2e-06 w=6e-06 

m1763 772 106 770 0 nenh l=2e-06 w=8e-06 

m1764 765 773 769 0 nenh l=2e-06 w=6e-06 

m1765 769 766 772 0 nenh l=2e-06 w=6e-06 

m1766 774 771 775 0 nenh l=2e-06 w=8e-06 

m1767 775 106 776 0 nenh l=2e-06 w=4e-06 

m1768 776 768 774 0 nenh l=2e-06 w=8e-06 

m1769 774 773 777 0 nenh l=2e-06 w=1e-05 

m1770 0 775 433 0 nenh l=2e-06 w=6e-06 

m1771 3 329 775 3 penh l=2e-06 w=1e-05 

m1772 775 433 3 3 penh l=8e-06 w=4e-06 

m1773 3 775 433 3 penh l=2e-06 w=1.6e-05 

m1774 3 778 757 3 penh l=2e-06 w=1.6e-05 

m1775 3 329 778 3 penh l=2e-06 w=1e-05 

m1776 778 757 3 3 penh l=8e-06 w=4e-06 

m1777 757 778 0 0 nenh l=2e-06 w=6e-06 

m1778 0 329 777 0 nenh l=2e-06 w=1.4e-05 

m1779 777 766 779 0 nenh l=2e-06 w=1.2e-05 

m1780 779 771 776 0 nenh l=2e-06 w=6e-06 

m1781 776 111 778 0 nenh l=2e-06 w=4e-06 

m1782 778 768 779 0 nenh l=2e-06 w=6e-06 

m1783 780 773 781 0 nenh l=2e-06 w=8e-06 

m1784 781 768 782 0 nenh l=2e-06 w=6e-06 

m1785 782 766 780 0 nenh l=2e-06 w=8e-06 

m1786 780 111 783 0 nenh l=2e-06 w=1e-05 

m1787 0 781 507 0 nenh l=2e-06 w=6e-06 

m1788 3 329 781 3 penh l=2e-06 w=1e-05 

m1789 781 507 3 3 penh l=8e-06 w=4e-06 

m1790 3 781 507 3 penh l=2e-06 w=1.6e-05 

m1791 3 784 512 3 penh l=2e-06 w=1.6e-05 

m1792 3 329 784 3 penh l=2e-06 w=1e-05 

m1793 784 512 3 3 penh l=8e-06 w=4e-06 

m1794 512 784 0 0 nenh l=2e-06 w=6e-06 

m1795 0 329 783 0 nenh l=2e-06 w=1.4e-05 

m1796 783 106 785 0 nenh l=2e-06 w=1e-05 

m1797 785 766 781 0 nenh l=2e-06 w=8e-06 

m1798 781 771 786 0 nenh l=2e-06 w=6e-06 

m1799 786 773 785 0 nenh l=2e-06 w=8e-06 

m1800 782 771 784 0 nenh l=2e-06 w=6e-06 

m1801 784 768 786 0 nenh l=2e-06 w=6e-06 

m1802 787 771 788 0 nenh l=2e-06 w=8e-06 

m1803 788 111 789 0 nenh l=2e-06 w=6e-06 

m1804 789 768 787 0 nenh l=2e-06 w=8e-06 

m1805 787 766 790 0 nenh l=2e-06 w=1e-05 

m1806 0 788 488 0 nenh l=2e-06 w=6e-06 

m1807 488 788 3 3 penh l=2e-06 w=1.6e-05 

m1808 3 488 788 3 penh l=8e-06 w=4e-06 

m1809 788 329 3 3 penh l=2e-06 w=1e-05 

m1810 3 791 499 3 penh l=2e-06 w=1.6e-05 

m1811 3 499 791 3 penh l=8e-06 w=4e-06 

m1812 791 329 3 3 penh l=2e-06 w=1e-05 

m1813 499 791 0 0 nenh l=2e-06 w=6e-06 

m1814 0 329 790 0 nenh l=2e-06 w=1.4e-05 

m1815 790 773 792 0 nenh l=2e-06 w=1e-05 

m1816 792 768 788 0 nenh l=2e-06 w=8e-06 

m1817 788 106 793 0 nenh l=2e-06 w=6e-06 

m1818 793 771 792 0 nenh l=2e-06 w=8e-06 

m1819 789 106 791 0 nenh l=2e-06 w=6e-06 

m1820 791 111 793 0 nenh l=2e-06 w=6e-06 

m1821 794 327 795 3 penh l=2e-06 w=5e-06 

m1822 795 329 796 3 penh l=2e-06 w=5e-06 

m1823 796 797 3 3 penh l=2e-06 w=5e-06 

m1824 3 795 797 3 penh l=2e-06 w=6e-06 

m1825 797 28 3 3 penh l=2e-06 w=6e-06 

m1826 3 797 305 3 penh l=2e-06 w=2.5e-05 

m1827 794 329 795 0 nenh l=2e-06 w=5e-06 

m1828 795 327 798 0 nenh l=2e-06 w=5e-06 

m1829 798 797 0 0 nenh l=2e-06 w=5e-06 

m1830 0 795 799 0 nenh l=2e-06 w=1.3e-05 

m1831 799 28 797 0 nenh l=2e-06 w=1.2e-05 

m1832 0 797 305 0 nenh l=2e-06 w=1.4e-05 

m1833 800 86 801 0 nenh l=2e-06 w=8e-06 

m1834 801 803 802 0 nenh l=2e-06 w=6e-06 

m1835 802 91 800 0 nenh l=2e-06 w=8e-06 

m1836 800 805 804 0 nenh l=2e-06 w=1e-05 

m1837 0 801 526 0 nenh l=2e-06 w=6e-06 

m1838 526 801 3 3 penh l=2e-06 w=1.6e-05 

m1839 3 526 801 3 penh l=8e-06 w=4e-06 

m1840 801 329 3 3 penh l=2e-06 w=1e-05 

m1841 3 806 534 3 penh l=2e-06 w=1.6e-05 

m1842 3 534 806 3 penh l=8e-06 w=4e-06 

m1843 806 329 3 3 penh l=2e-06 w=1e-05 

m1844 534 806 0 0 nenh l=2e-06 w=6e-06 

m1845 0 329 804 0 nenh l=2e-06 w=1.4e-05 

m1846 804 808 807 0 nenh l=2e-06 w=1e-05 

m1847 807 91 801 0 nenh l=2e-06 w=8e-06 

m1848 801 810 809 0 nenh l=2e-06 w=6e-06 

m1849 809 86 807 0 nenh l=2e-06 w=8e-06 

m1850 802 810 806 0 nenh l=2e-06 w=6e-06 

m1851 806 803 809 0 nenh l=2e-06 w=6e-06 

m1852 811 808 812 0 nenh l=2e-06 w=8e-06 

m1853 812 86 813 0 nenh l=2e-06 w=4e-06 

m1854 813 805 811 0 nenh l=2e-06 w=8e-06 

m1855 811 810 814 0 nenh l=2e-06 w=1e-05 

m1856 0 812 436 0 nenh l=2e-06 w=6e-06 

m1857 3 329 812 3 penh l=2e-06 w=1e-05 

m1858 812 436 3 3 penh l=8e-06 w=4e-06 

m1859 3 812 436 3 penh l=2e-06 w=1.6e-05 

m1860 3 815 794 3 penh l=2e-06 w=1.6e-05 

m1861 3 329 815 3 penh l=2e-06 w=1e-05 

m1862 815 794 3 3 penh l=8e-06 w=4e-06 

m1863 794 815 0 0 nenh l=2e-06 w=6e-06 

m1864 0 329 814 0 nenh l=2e-06 w=1.4e-05 

m1865 814 803 816 0 nenh l=2e-06 w=1.2e-05 

m1866 816 808 813 0 nenh l=2e-06 w=6e-06 

m1867 813 91 815 0 nenh l=2e-06 w=4e-06 

m1868 815 805 816 0 nenh l=2e-06 w=6e-06 

m1869 817 810 818 0 nenh l=2e-06 w=8e-06 

m1870 818 805 819 0 nenh l=2e-06 w=6e-06 

m1871 819 803 817 0 nenh l=2e-06 w=8e-06 

m1872 817 91 820 0 nenh l=2e-06 w=1e-05 

m1873 0 818 509 0 nenh l=2e-06 w=6e-06 

m1874 3 329 818 3 penh l=2e-06 w=1e-05 

m1875 818 509 3 3 penh l=8e-06 w=4e-06 

m1876 3 818 509 3 penh l=2e-06 w=1.6e-05 

m1877 3 821 517 3 penh l=2e-06 w=1.6e-05 

m1878 3 329 821 3 penh l=2e-06 w=1e-05 

m1879 821 517 3 3 penh l=8e-06 w=4e-06 

m1880 517 821 0 0 nenh l=2e-06 w=6e-06 

m1881 0 329 820 0 nenh l=2e-06 w=1.4e-05 

m1882 820 86 822 0 nenh l=2e-06 w=1e-05 

m1883 822 803 818 0 nenh l=2e-06 w=8e-06 

m1884 818 808 823 0 nenh l=2e-06 w=6e-06 

m1885 823 810 822 0 nenh l=2e-06 w=8e-06 

m1886 819 808 821 0 nenh l=2e-06 w=6e-06 

m1887 821 805 823 0 nenh l=2e-06 w=6e-06 

m1888 824 808 825 0 nenh l=2e-06 w=8e-06 

m1889 825 91 826 0 nenh l=2e-06 w=6e-06 

m1890 826 805 824 0 nenh l=2e-06 w=8e-06 

m1891 824 803 827 0 nenh l=2e-06 w=1e-05 

m1892 0 825 486 0 nenh l=2e-06 w=6e-06 

m1893 486 825 3 3 penh l=2e-06 w=1.6e-05 

m1894 3 486 825 3 penh l=8e-06 w=4e-06 

m1895 825 329 3 3 penh l=2e-06 w=1e-05 

m1896 3 828 498 3 penh l=2e-06 w=1.6e-05 

m1897 3 498 828 3 penh l=8e-06 w=4e-06 

m1898 828 329 3 3 penh l=2e-06 w=1e-05 

m1899 498 828 0 0 nenh l=2e-06 w=6e-06 

m1900 0 329 827 0 nenh l=2e-06 w=1.4e-05 

m1901 827 810 829 0 nenh l=2e-06 w=1e-05 

m1902 829 805 825 0 nenh l=2e-06 w=8e-06 

m1903 825 86 830 0 nenh l=2e-06 w=6e-06 

m1904 830 808 829 0 nenh l=2e-06 w=8e-06 

m1905 826 86 828 0 nenh l=2e-06 w=6e-06 

m1906 828 91 830 0 nenh l=2e-06 w=6e-06 

m1907 132 831 3 3 penh l=2e-06 w=6.2e-05 

m1908 3 832 831 3 penh l=2e-06 w=6.2e-05 

m1909 832 833 3 3 penh l=2e-06 w=2.9e-05 

m1910 3 834 833 3 penh l=4e-06 w=2.9e-05 

m1911 832 833 0 0 nenh l=2e-06 w=2.1e-05 

m1912 0 834 833 0 nenh l=4e-06 w=2.1e-05 

m1913 132 831 0 0 nenh l=2e-06 w=4.8e-05 

m1914 0 832 831 0 nenh l=2e-06 w=4.8e-05 

m1915 834 0 0 0 nenh l=4e-06 w=2.5e-05 

m1916 112 835 3 3 penh l=2e-06 w=6.2e-05 

m1917 3 836 835 3 penh l=2e-06 w=6.2e-05 

m1918 836 837 3 3 penh l=2e-06 w=2.9e-05 

m1919 3 838 837 3 penh l=4e-06 w=2.9e-05 

m1920 836 837 0 0 nenh l=2e-06 w=2.1e-05 

m1921 0 838 837 0 nenh l=4e-06 w=2.1e-05 

m1922 112 835 0 0 nenh l=2e-06 w=4.8e-05 

m1923 0 836 835 0 nenh l=2e-06 w=4.8e-05 

m1924 838 0 0 0 nenh l=4e-06 w=2.5e-05 

m1925 3 840 839 3 penh l=2e-06 w=9.7e-05 

m1926 839 840 3 3 penh l=2e-06 w=9.5e-05 

m1927 3 840 839 3 penh l=2e-06 w=9.5e-05 

m1928 839 840 3 3 penh l=2e-06 w=9.6e-05 

m1929 3 840 839 3 penh l=2e-06 w=9.6e-05 

m1930 839 840 3 3 penh l=2e-06 w=9.5e-05 

m1931 3 840 839 3 penh l=2e-06 w=9.5e-05 

m1932 839 840 3 3 penh l=2e-06 w=9.6e-05 

m1933 3 841 840 3 penh l=2e-06 w=5.3e-05 

m1934 840 841 3 3 penh l=2e-06 w=5.3e-05 

m1935 3 842 841 3 penh l=2e-06 w=4.9e-05 

m1936 842 292 3 3 penh l=2e-06 w=2.3e-05 

m1937 3 841 840 3 penh l=2e-06 w=4.8e-05 

m1938 840 841 3 3 penh l=2e-06 w=4.8e-05 

m1939 3 292 843 3 penh l=2e-06 w=2.2e-05 

m1940 844 845 3 3 penh l=2e-06 w=5e-05 

m1941 3 843 845 3 penh l=2e-06 w=4.7e-05 

m1942 844 845 3 3 penh l=2e-06 w=4.8e-05 

m1943 3 845 844 3 penh l=2e-06 w=4.8e-05 

m1944 0 844 839 0 nenh l=2e-06 w=4.6e-05 

m1945 839 844 0 0 nenh l=2e-06 w=4.8e-05 

m1946 0 844 839 0 nenh l=2e-06 w=4.6e-05 

m1947 839 844 0 0 nenh l=2e-06 w=4.8e-05 

m1948 0 844 839 0 nenh l=2e-06 w=4.8e-05 

m1949 839 844 0 0 nenh l=2e-06 w=4.8e-05 

m1950 0 844 839 0 nenh l=2e-06 w=4.8e-05 

m1951 839 844 0 0 nenh l=2e-06 w=4.6e-05 

m1952 0 845 844 0 nenh l=2e-06 w=6e-05 

m1953 844 845 0 0 nenh l=2e-06 w=6e-05 

m1954 845 843 0 0 nenh l=2e-06 w=5e-05 

m1955 0 841 840 0 nenh l=2e-06 w=3.5e-05 

m1956 840 841 0 0 nenh l=2e-06 w=3.4e-05 

m1957 0 292 843 0 nenh l=2e-06 w=2.4e-05 

m1958 0 841 840 0 nenh l=2e-06 w=2.5e-05 

m1959 840 841 0 0 nenh l=2e-06 w=2.5e-05 

m1960 0 842 841 0 nenh l=2e-06 w=1.6e-05 

m1961 842 292 0 0 nenh l=2e-06 w=2.3e-05 

m1962 3 847 846 3 penh l=2e-06 w=9.7e-05 

m1963 846 847 3 3 penh l=2e-06 w=9.5e-05 

m1964 3 847 846 3 penh l=2e-06 w=9.5e-05 

m1965 846 847 3 3 penh l=2e-06 w=9.6e-05 

m1966 3 847 846 3 penh l=2e-06 w=9.6e-05 

m1967 846 847 3 3 penh l=2e-06 w=9.5e-05 

m1968 3 847 846 3 penh l=2e-06 w=9.5e-05 

m1969 846 847 3 3 penh l=2e-06 w=9.6e-05 

m1970 3 848 847 3 penh l=2e-06 w=5.3e-05 

m1971 847 848 3 3 penh l=2e-06 w=5.3e-05 

m1972 3 849 848 3 penh l=2e-06 w=4.9e-05 

m1973 849 287 3 3 penh l=2e-06 w=2.3e-05 

m1974 3 848 847 3 penh l=2e-06 w=4.8e-05 

m1975 847 848 3 3 penh l=2e-06 w=4.8e-05 

m1976 3 287 850 3 penh l=2e-06 w=2.2e-05 

m1977 851 852 3 3 penh l=2e-06 w=5e-05 

m1978 3 850 852 3 penh l=2e-06 w=4.7e-05 

m1979 851 852 3 3 penh l=2e-06 w=4.8e-05 

m1980 3 852 851 3 penh l=2e-06 w=4.8e-05 

m1981 0 851 846 0 nenh l=2e-06 w=4.6e-05 

m1982 846 851 0 0 nenh l=2e-06 w=4.8e-05 

m1983 0 851 846 0 nenh l=2e-06 w=4.6e-05 

m1984 846 851 0 0 nenh l=2e-06 w=4.8e-05 

m1985 0 851 846 0 nenh l=2e-06 w=4.8e-05 

m1986 846 851 0 0 nenh l=2e-06 w=4.8e-05 

m1987 0 851 846 0 nenh l=2e-06 w=4.8e-05 

m1988 846 851 0 0 nenh l=2e-06 w=4.6e-05 

m1989 0 852 851 0 nenh l=2e-06 w=6e-05 

m1990 851 852 0 0 nenh l=2e-06 w=6e-05 

m1991 852 850 0 0 nenh l=2e-06 w=5e-05 

m1992 0 848 847 0 nenh l=2e-06 w=3.5e-05 

m1993 847 848 0 0 nenh l=2e-06 w=3.4e-05 

m1994 0 287 850 0 nenh l=2e-06 w=2.4e-05 

m1995 0 848 847 0 nenh l=2e-06 w=2.5e-05 

m1996 847 848 0 0 nenh l=2e-06 w=2.5e-05 

m1997 0 849 848 0 nenh l=2e-06 w=1.6e-05 

m1998 849 287 0 0 nenh l=2e-06 w=2.3e-05 

m1999 853 327 854 3 penh l=2e-06 w=5e-06 

m2000 854 329 855 3 penh l=2e-06 w=5e-06 

m2001 855 856 3 3 penh l=2e-06 w=5e-06 

m2002 3 854 856 3 penh l=2e-06 w=6e-06 

m2003 856 857 3 3 penh l=2e-06 w=6e-06 

m2004 3 856 274 3 penh l=2e-06 w=2.5e-05 

m2005 853 329 854 0 nenh l=2e-06 w=5e-06 

m2006 854 327 858 0 nenh l=2e-06 w=5e-06 

m2007 858 856 0 0 nenh l=2e-06 w=5e-06 

m2008 0 854 859 0 nenh l=2e-06 w=1.3e-05 

m2009 859 857 856 0 nenh l=2e-06 w=1.2e-05 

m2010 0 856 274 0 nenh l=2e-06 w=1.4e-05 

m2011 860 223 861 0 nenh l=2e-06 w=8e-06 

m2012 861 544 862 0 nenh l=2e-06 w=6e-06 

m2013 862 228 860 0 nenh l=2e-06 w=8e-06 

m2014 860 546 863 0 nenh l=2e-06 w=1e-05 

m2015 0 861 864 0 nenh l=2e-06 w=6e-06 

m2016 864 861 3 3 penh l=2e-06 w=1.6e-05 

m2017 3 864 861 3 penh l=8e-06 w=4e-06 

m2018 861 329 3 3 penh l=2e-06 w=1e-05 

m2019 3 866 865 3 penh l=2e-06 w=1.6e-05 

m2020 3 865 866 3 penh l=8e-06 w=4e-06 

m2021 866 329 3 3 penh l=2e-06 w=1e-05 

m2022 865 866 0 0 nenh l=2e-06 w=6e-06 

m2023 0 329 863 0 nenh l=2e-06 w=1.4e-05 

m2024 863 549 867 0 nenh l=2e-06 w=1e-05 

m2025 867 228 861 0 nenh l=2e-06 w=8e-06 

m2026 861 551 868 0 nenh l=2e-06 w=6e-06 

m2027 868 223 867 0 nenh l=2e-06 w=8e-06 

m2028 862 551 866 0 nenh l=2e-06 w=6e-06 

m2029 866 544 868 0 nenh l=2e-06 w=6e-06 

m2030 869 549 870 0 nenh l=2e-06 w=8e-06 

m2031 870 223 871 0 nenh l=2e-06 w=4e-06 

m2032 871 546 869 0 nenh l=2e-06 w=8e-06 

m2033 869 551 872 0 nenh l=2e-06 w=1e-05 

m2034 0 870 873 0 nenh l=2e-06 w=6e-06 

m2035 3 329 870 3 penh l=2e-06 w=1e-05 

m2036 870 873 3 3 penh l=8e-06 w=4e-06 

m2037 3 870 873 3 penh l=2e-06 w=1.6e-05 

m2038 3 874 853 3 penh l=2e-06 w=1.6e-05 

m2039 3 329 874 3 penh l=2e-06 w=1e-05 

m2040 874 853 3 3 penh l=8e-06 w=4e-06 

m2041 853 874 0 0 nenh l=2e-06 w=6e-06 

m2042 0 329 872 0 nenh l=2e-06 w=1.4e-05 

m2043 872 544 875 0 nenh l=2e-06 w=1.2e-05 

m2044 875 549 871 0 nenh l=2e-06 w=6e-06 

m2045 871 228 874 0 nenh l=2e-06 w=4e-06 

m2046 874 546 875 0 nenh l=2e-06 w=6e-06 

m2047 876 551 877 0 nenh l=2e-06 w=8e-06 

m2048 877 546 878 0 nenh l=2e-06 w=6e-06 

m2049 878 544 876 0 nenh l=2e-06 w=8e-06 

m2050 876 228 879 0 nenh l=2e-06 w=1e-05 

m2051 0 877 880 0 nenh l=2e-06 w=6e-06 

m2052 3 329 877 3 penh l=2e-06 w=1e-05 

m2053 877 880 3 3 penh l=8e-06 w=4e-06 

m2054 3 877 880 3 penh l=2e-06 w=1.6e-05 

m2055 3 882 881 3 penh l=2e-06 w=1.6e-05 

m2056 3 329 882 3 penh l=2e-06 w=1e-05 

m2057 882 881 3 3 penh l=8e-06 w=4e-06 

m2058 881 882 0 0 nenh l=2e-06 w=6e-06 

m2059 0 329 879 0 nenh l=2e-06 w=1.4e-05 

m2060 879 223 883 0 nenh l=2e-06 w=1e-05 

m2061 883 544 877 0 nenh l=2e-06 w=8e-06 

m2062 877 549 884 0 nenh l=2e-06 w=6e-06 

m2063 884 551 883 0 nenh l=2e-06 w=8e-06 

m2064 878 549 882 0 nenh l=2e-06 w=6e-06 

m2065 882 546 884 0 nenh l=2e-06 w=6e-06 

m2066 885 549 886 0 nenh l=2e-06 w=8e-06 

m2067 886 228 887 0 nenh l=2e-06 w=6e-06 

m2068 887 546 885 0 nenh l=2e-06 w=8e-06 

m2069 885 544 888 0 nenh l=2e-06 w=1e-05 

m2070 0 886 889 0 nenh l=2e-06 w=6e-06 

m2071 889 886 3 3 penh l=2e-06 w=1.6e-05 

m2072 3 889 886 3 penh l=8e-06 w=4e-06 

m2073 886 329 3 3 penh l=2e-06 w=1e-05 

m2074 3 891 890 3 penh l=2e-06 w=1.6e-05 

m2075 3 890 891 3 penh l=8e-06 w=4e-06 

m2076 891 329 3 3 penh l=2e-06 w=1e-05 

m2077 890 891 0 0 nenh l=2e-06 w=6e-06 

m2078 0 329 888 0 nenh l=2e-06 w=1.4e-05 

m2079 888 551 892 0 nenh l=2e-06 w=1e-05 

m2080 892 546 886 0 nenh l=2e-06 w=8e-06 

m2081 886 223 893 0 nenh l=2e-06 w=6e-06 

m2082 893 549 892 0 nenh l=2e-06 w=8e-06 

m2083 887 223 891 0 nenh l=2e-06 w=6e-06 

m2084 891 228 893 0 nenh l=2e-06 w=6e-06 

m2085 894 327 895 3 penh l=2e-06 w=5e-06 

m2086 895 329 896 3 penh l=2e-06 w=5e-06 

m2087 896 897 3 3 penh l=2e-06 w=5e-06 

m2088 3 895 897 3 penh l=2e-06 w=6e-06 

m2089 897 857 3 3 penh l=2e-06 w=6e-06 

m2090 3 897 280 3 penh l=2e-06 w=2.5e-05 

m2091 894 329 895 0 nenh l=2e-06 w=5e-06 

m2092 895 327 898 0 nenh l=2e-06 w=5e-06 

m2093 898 897 0 0 nenh l=2e-06 w=5e-06 

m2094 0 895 899 0 nenh l=2e-06 w=1.3e-05 

m2095 899 857 897 0 nenh l=2e-06 w=1.2e-05 

m2096 0 897 280 0 nenh l=2e-06 w=1.4e-05 

m2097 900 204 901 0 nenh l=2e-06 w=8e-06 

m2098 901 581 902 0 nenh l=2e-06 w=6e-06 

m2099 902 209 900 0 nenh l=2e-06 w=8e-06 

m2100 900 583 903 0 nenh l=2e-06 w=1e-05 

m2101 0 901 904 0 nenh l=2e-06 w=6e-06 

m2102 904 901 3 3 penh l=2e-06 w=1.6e-05 

m2103 3 904 901 3 penh l=8e-06 w=4e-06 

m2104 901 329 3 3 penh l=2e-06 w=1e-05 

m2105 3 906 905 3 penh l=2e-06 w=1.6e-05 

m2106 3 905 906 3 penh l=8e-06 w=4e-06 

m2107 906 329 3 3 penh l=2e-06 w=1e-05 

m2108 905 906 0 0 nenh l=2e-06 w=6e-06 

m2109 0 329 903 0 nenh l=2e-06 w=1.4e-05 

m2110 903 586 907 0 nenh l=2e-06 w=1e-05 

m2111 907 209 901 0 nenh l=2e-06 w=8e-06 

m2112 901 588 908 0 nenh l=2e-06 w=6e-06 

m2113 908 204 907 0 nenh l=2e-06 w=8e-06 

m2114 902 588 906 0 nenh l=2e-06 w=6e-06 

m2115 906 581 908 0 nenh l=2e-06 w=6e-06 

m2116 909 586 910 0 nenh l=2e-06 w=8e-06 

m2117 910 204 911 0 nenh l=2e-06 w=4e-06 

m2118 911 583 909 0 nenh l=2e-06 w=8e-06 

m2119 909 588 912 0 nenh l=2e-06 w=1e-05 

m2120 0 910 913 0 nenh l=2e-06 w=6e-06 

m2121 3 329 910 3 penh l=2e-06 w=1e-05 

m2122 910 913 3 3 penh l=8e-06 w=4e-06 

m2123 3 910 913 3 penh l=2e-06 w=1.6e-05 

m2124 3 914 894 3 penh l=2e-06 w=1.6e-05 

m2125 3 329 914 3 penh l=2e-06 w=1e-05 

m2126 914 894 3 3 penh l=8e-06 w=4e-06 

m2127 894 914 0 0 nenh l=2e-06 w=6e-06 

m2128 0 329 912 0 nenh l=2e-06 w=1.4e-05 

m2129 912 581 915 0 nenh l=2e-06 w=1.2e-05 

m2130 915 586 911 0 nenh l=2e-06 w=6e-06 

m2131 911 209 914 0 nenh l=2e-06 w=4e-06 

m2132 914 583 915 0 nenh l=2e-06 w=6e-06 

m2133 916 588 917 0 nenh l=2e-06 w=8e-06 

m2134 917 583 918 0 nenh l=2e-06 w=6e-06 

m2135 918 581 916 0 nenh l=2e-06 w=8e-06 

m2136 916 209 919 0 nenh l=2e-06 w=1e-05 

m2137 0 917 920 0 nenh l=2e-06 w=6e-06 

m2138 3 329 917 3 penh l=2e-06 w=1e-05 

m2139 917 920 3 3 penh l=8e-06 w=4e-06 

m2140 3 917 920 3 penh l=2e-06 w=1.6e-05 

m2141 3 922 921 3 penh l=2e-06 w=1.6e-05 

m2142 3 329 922 3 penh l=2e-06 w=1e-05 

m2143 922 921 3 3 penh l=8e-06 w=4e-06 

m2144 921 922 0 0 nenh l=2e-06 w=6e-06 

m2145 0 329 919 0 nenh l=2e-06 w=1.4e-05 

m2146 919 204 923 0 nenh l=2e-06 w=1e-05 

m2147 923 581 917 0 nenh l=2e-06 w=8e-06 

m2148 917 586 924 0 nenh l=2e-06 w=6e-06 

m2149 924 588 923 0 nenh l=2e-06 w=8e-06 

m2150 918 586 922 0 nenh l=2e-06 w=6e-06 

m2151 922 583 924 0 nenh l=2e-06 w=6e-06 

m2152 925 586 926 0 nenh l=2e-06 w=8e-06 

m2153 926 209 927 0 nenh l=2e-06 w=6e-06 

m2154 927 583 925 0 nenh l=2e-06 w=8e-06 

m2155 925 581 928 0 nenh l=2e-06 w=1e-05 

m2156 0 926 929 0 nenh l=2e-06 w=6e-06 

m2157 929 926 3 3 penh l=2e-06 w=1.6e-05 

m2158 3 929 926 3 penh l=8e-06 w=4e-06 

m2159 926 329 3 3 penh l=2e-06 w=1e-05 

m2160 3 931 930 3 penh l=2e-06 w=1.6e-05 

m2161 3 930 931 3 penh l=8e-06 w=4e-06 

m2162 931 329 3 3 penh l=2e-06 w=1e-05 

m2163 930 931 0 0 nenh l=2e-06 w=6e-06 

m2164 0 329 928 0 nenh l=2e-06 w=1.4e-05 

m2165 928 588 932 0 nenh l=2e-06 w=1e-05 

m2166 932 583 926 0 nenh l=2e-06 w=8e-06 

m2167 926 204 933 0 nenh l=2e-06 w=6e-06 

m2168 933 586 932 0 nenh l=2e-06 w=8e-06 

m2169 927 204 931 0 nenh l=2e-06 w=6e-06 

m2170 931 209 933 0 nenh l=2e-06 w=6e-06 

m2171 934 327 935 3 penh l=2e-06 w=5e-06 

m2172 935 329 936 3 penh l=2e-06 w=5e-06 

m2173 936 937 3 3 penh l=2e-06 w=5e-06 

m2174 3 935 937 3 penh l=2e-06 w=6e-06 

m2175 937 857 3 3 penh l=2e-06 w=6e-06 

m2176 3 937 285 3 penh l=2e-06 w=2.5e-05 

m2177 934 329 935 0 nenh l=2e-06 w=5e-06 

m2178 935 327 938 0 nenh l=2e-06 w=5e-06 

m2179 938 937 0 0 nenh l=2e-06 w=5e-06 

m2180 0 935 939 0 nenh l=2e-06 w=1.3e-05 

m2181 939 857 937 0 nenh l=2e-06 w=1.2e-05 

m2182 0 937 285 0 nenh l=2e-06 w=1.4e-05 

m2183 940 185 941 0 nenh l=2e-06 w=8e-06 

m2184 941 618 942 0 nenh l=2e-06 w=6e-06 

m2185 942 190 940 0 nenh l=2e-06 w=8e-06 

m2186 940 620 943 0 nenh l=2e-06 w=1e-05 

m2187 0 941 944 0 nenh l=2e-06 w=6e-06 

m2188 944 941 3 3 penh l=2e-06 w=1.6e-05 

m2189 3 944 941 3 penh l=8e-06 w=4e-06 

m2190 941 329 3 3 penh l=2e-06 w=1e-05 

m2191 3 946 945 3 penh l=2e-06 w=1.6e-05 

m2192 3 945 946 3 penh l=8e-06 w=4e-06 

m2193 946 329 3 3 penh l=2e-06 w=1e-05 

m2194 945 946 0 0 nenh l=2e-06 w=6e-06 

m2195 0 329 943 0 nenh l=2e-06 w=1.4e-05 

m2196 943 623 947 0 nenh l=2e-06 w=1e-05 

m2197 947 190 941 0 nenh l=2e-06 w=8e-06 

m2198 941 625 948 0 nenh l=2e-06 w=6e-06 

m2199 948 185 947 0 nenh l=2e-06 w=8e-06 

m2200 942 625 946 0 nenh l=2e-06 w=6e-06 

m2201 946 618 948 0 nenh l=2e-06 w=6e-06 

m2202 949 623 950 0 nenh l=2e-06 w=8e-06 

m2203 950 185 951 0 nenh l=2e-06 w=4e-06 

m2204 951 620 949 0 nenh l=2e-06 w=8e-06 

m2205 949 625 952 0 nenh l=2e-06 w=1e-05 

m2206 0 950 953 0 nenh l=2e-06 w=6e-06 

m2207 3 329 950 3 penh l=2e-06 w=1e-05 

m2208 950 953 3 3 penh l=8e-06 w=4e-06 

m2209 3 950 953 3 penh l=2e-06 w=1.6e-05 

m2210 3 954 934 3 penh l=2e-06 w=1.6e-05 

m2211 3 329 954 3 penh l=2e-06 w=1e-05 

m2212 954 934 3 3 penh l=8e-06 w=4e-06 

m2213 934 954 0 0 nenh l=2e-06 w=6e-06 

m2214 0 329 952 0 nenh l=2e-06 w=1.4e-05 

m2215 952 618 955 0 nenh l=2e-06 w=1.2e-05 

m2216 955 623 951 0 nenh l=2e-06 w=6e-06 

m2217 951 190 954 0 nenh l=2e-06 w=4e-06 

m2218 954 620 955 0 nenh l=2e-06 w=6e-06 

m2219 956 625 957 0 nenh l=2e-06 w=8e-06 

m2220 957 620 958 0 nenh l=2e-06 w=6e-06 

m2221 958 618 956 0 nenh l=2e-06 w=8e-06 

m2222 956 190 959 0 nenh l=2e-06 w=1e-05 

m2223 0 957 960 0 nenh l=2e-06 w=6e-06 

m2224 3 329 957 3 penh l=2e-06 w=1e-05 

m2225 957 960 3 3 penh l=8e-06 w=4e-06 

m2226 3 957 960 3 penh l=2e-06 w=1.6e-05 

m2227 3 962 961 3 penh l=2e-06 w=1.6e-05 

m2228 3 329 962 3 penh l=2e-06 w=1e-05 

m2229 962 961 3 3 penh l=8e-06 w=4e-06 

m2230 961 962 0 0 nenh l=2e-06 w=6e-06 

m2231 0 329 959 0 nenh l=2e-06 w=1.4e-05 

m2232 959 185 963 0 nenh l=2e-06 w=1e-05 

m2233 963 618 957 0 nenh l=2e-06 w=8e-06 

m2234 957 623 964 0 nenh l=2e-06 w=6e-06 

m2235 964 625 963 0 nenh l=2e-06 w=8e-06 

m2236 958 623 962 0 nenh l=2e-06 w=6e-06 

m2237 962 620 964 0 nenh l=2e-06 w=6e-06 

m2238 965 623 966 0 nenh l=2e-06 w=8e-06 

m2239 966 190 967 0 nenh l=2e-06 w=6e-06 

m2240 967 620 965 0 nenh l=2e-06 w=8e-06 

m2241 965 618 968 0 nenh l=2e-06 w=1e-05 

m2242 0 966 969 0 nenh l=2e-06 w=6e-06 

m2243 969 966 3 3 penh l=2e-06 w=1.6e-05 

m2244 3 969 966 3 penh l=8e-06 w=4e-06 

m2245 966 329 3 3 penh l=2e-06 w=1e-05 

m2246 3 971 970 3 penh l=2e-06 w=1.6e-05 

m2247 3 970 971 3 penh l=8e-06 w=4e-06 

m2248 971 329 3 3 penh l=2e-06 w=1e-05 

m2249 970 971 0 0 nenh l=2e-06 w=6e-06 

m2250 0 329 968 0 nenh l=2e-06 w=1.4e-05 

m2251 968 625 972 0 nenh l=2e-06 w=1e-05 

m2252 972 620 966 0 nenh l=2e-06 w=8e-06 

m2253 966 185 973 0 nenh l=2e-06 w=6e-06 

m2254 973 623 972 0 nenh l=2e-06 w=8e-06 

m2255 967 185 971 0 nenh l=2e-06 w=6e-06 

m2256 971 190 973 0 nenh l=2e-06 w=6e-06 

m2257 974 327 975 3 penh l=2e-06 w=5e-06 

m2258 975 329 976 3 penh l=2e-06 w=5e-06 

m2259 976 977 3 3 penh l=2e-06 w=5e-06 

m2260 3 975 977 3 penh l=2e-06 w=6e-06 

m2261 977 857 3 3 penh l=2e-06 w=6e-06 

m2262 3 977 290 3 penh l=2e-06 w=2.5e-05 

m2263 974 329 975 0 nenh l=2e-06 w=5e-06 

m2264 975 327 978 0 nenh l=2e-06 w=5e-06 

m2265 978 977 0 0 nenh l=2e-06 w=5e-06 

m2266 0 975 979 0 nenh l=2e-06 w=1.3e-05 

m2267 979 857 977 0 nenh l=2e-06 w=1.2e-05 

m2268 0 977 290 0 nenh l=2e-06 w=1.4e-05 

m2269 980 166 981 0 nenh l=2e-06 w=8e-06 

m2270 981 655 982 0 nenh l=2e-06 w=6e-06 

m2271 982 171 980 0 nenh l=2e-06 w=8e-06 

m2272 980 657 983 0 nenh l=2e-06 w=1e-05 

m2273 0 981 984 0 nenh l=2e-06 w=6e-06 

m2274 984 981 3 3 penh l=2e-06 w=1.6e-05 

m2275 3 984 981 3 penh l=8e-06 w=4e-06 

m2276 981 329 3 3 penh l=2e-06 w=1e-05 

m2277 3 986 985 3 penh l=2e-06 w=1.6e-05 

m2278 3 985 986 3 penh l=8e-06 w=4e-06 

m2279 986 329 3 3 penh l=2e-06 w=1e-05 

m2280 985 986 0 0 nenh l=2e-06 w=6e-06 

m2281 0 329 983 0 nenh l=2e-06 w=1.4e-05 

m2282 983 660 987 0 nenh l=2e-06 w=1e-05 

m2283 987 171 981 0 nenh l=2e-06 w=8e-06 

m2284 981 662 988 0 nenh l=2e-06 w=6e-06 

m2285 988 166 987 0 nenh l=2e-06 w=8e-06 

m2286 982 662 986 0 nenh l=2e-06 w=6e-06 

m2287 986 655 988 0 nenh l=2e-06 w=6e-06 

m2288 989 660 990 0 nenh l=2e-06 w=8e-06 

m2289 990 166 991 0 nenh l=2e-06 w=4e-06 

m2290 991 657 989 0 nenh l=2e-06 w=8e-06 

m2291 989 662 992 0 nenh l=2e-06 w=1e-05 

m2292 0 990 993 0 nenh l=2e-06 w=6e-06 

m2293 3 329 990 3 penh l=2e-06 w=1e-05 

m2294 990 993 3 3 penh l=8e-06 w=4e-06 

m2295 3 990 993 3 penh l=2e-06 w=1.6e-05 

m2296 3 994 974 3 penh l=2e-06 w=1.6e-05 

m2297 3 329 994 3 penh l=2e-06 w=1e-05 

m2298 994 974 3 3 penh l=8e-06 w=4e-06 

m2299 974 994 0 0 nenh l=2e-06 w=6e-06 

m2300 0 329 992 0 nenh l=2e-06 w=1.4e-05 

m2301 992 655 995 0 nenh l=2e-06 w=1.2e-05 

m2302 995 660 991 0 nenh l=2e-06 w=6e-06 

m2303 991 171 994 0 nenh l=2e-06 w=4e-06 

m2304 994 657 995 0 nenh l=2e-06 w=6e-06 

m2305 996 662 997 0 nenh l=2e-06 w=8e-06 

m2306 997 657 998 0 nenh l=2e-06 w=6e-06 

m2307 998 655 996 0 nenh l=2e-06 w=8e-06 

m2308 996 171 999 0 nenh l=2e-06 w=1e-05 

m2309 0 997 1000 0 nenh l=2e-06 w=6e-06 

m2310 3 329 997 3 penh l=2e-06 w=1e-05 

m2311 997 1000 3 3 penh l=8e-06 w=4e-06 

m2312 3 997 1000 3 penh l=2e-06 w=1.6e-05 

m2313 3 1002 1001 3 penh l=2e-06 w=1.6e-05 

m2314 3 329 1002 3 penh l=2e-06 w=1e-05 

m2315 1002 1001 3 3 penh l=8e-06 w=4e-06 

m2316 1001 1002 0 0 nenh l=2e-06 w=6e-06 

m2317 0 329 999 0 nenh l=2e-06 w=1.4e-05 

m2318 999 166 1003 0 nenh l=2e-06 w=1e-05 

m2319 1003 655 997 0 nenh l=2e-06 w=8e-06 

m2320 997 660 1004 0 nenh l=2e-06 w=6e-06 

m2321 1004 662 1003 0 nenh l=2e-06 w=8e-06 

m2322 998 660 1002 0 nenh l=2e-06 w=6e-06 

m2323 1002 657 1004 0 nenh l=2e-06 w=6e-06 

m2324 1005 660 1006 0 nenh l=2e-06 w=8e-06 

m2325 1006 171 1007 0 nenh l=2e-06 w=6e-06 

m2326 1007 657 1005 0 nenh l=2e-06 w=8e-06 

m2327 1005 655 1008 0 nenh l=2e-06 w=1e-05 

m2328 0 1006 1009 0 nenh l=2e-06 w=6e-06 

m2329 1009 1006 3 3 penh l=2e-06 w=1.6e-05 

m2330 3 1009 1006 3 penh l=8e-06 w=4e-06 

m2331 1006 329 3 3 penh l=2e-06 w=1e-05 

m2332 3 1011 1010 3 penh l=2e-06 w=1.6e-05 

m2333 3 1010 1011 3 penh l=8e-06 w=4e-06 

m2334 1011 329 3 3 penh l=2e-06 w=1e-05 

m2335 1010 1011 0 0 nenh l=2e-06 w=6e-06 

m2336 0 329 1008 0 nenh l=2e-06 w=1.4e-05 

m2337 1008 662 1012 0 nenh l=2e-06 w=1e-05 

m2338 1012 657 1006 0 nenh l=2e-06 w=8e-06 

m2339 1006 166 1013 0 nenh l=2e-06 w=6e-06 

m2340 1013 660 1012 0 nenh l=2e-06 w=8e-06 

m2341 1007 166 1011 0 nenh l=2e-06 w=6e-06 

m2342 1011 171 1013 0 nenh l=2e-06 w=6e-06 

m2343 1014 327 1015 3 penh l=2e-06 w=5e-06 

m2344 1015 329 1016 3 penh l=2e-06 w=5e-06 

m2345 1016 1017 3 3 penh l=2e-06 w=5e-06 

m2346 3 1015 1017 3 penh l=2e-06 w=6e-06 

m2347 1017 857 3 3 penh l=2e-06 w=6e-06 

m2348 3 1017 295 3 penh l=2e-06 w=2.5e-05 

m2349 1014 329 1015 0 nenh l=2e-06 w=5e-06 

m2350 1015 327 1018 0 nenh l=2e-06 w=5e-06 

m2351 1018 1017 0 0 nenh l=2e-06 w=5e-06 

m2352 0 1015 1019 0 nenh l=2e-06 w=1.3e-05 

m2353 1019 857 1017 0 nenh l=2e-06 w=1.2e-05 

m2354 0 1017 295 0 nenh l=2e-06 w=1.4e-05 

m2355 1020 146 1021 0 nenh l=2e-06 w=8e-06 

m2356 1021 692 1022 0 nenh l=2e-06 w=6e-06 

m2357 1022 151 1020 0 nenh l=2e-06 w=8e-06 

m2358 1020 694 1023 0 nenh l=2e-06 w=1e-05 

m2359 0 1021 1024 0 nenh l=2e-06 w=6e-06 

m2360 1024 1021 3 3 penh l=2e-06 w=1.6e-05 

m2361 3 1024 1021 3 penh l=8e-06 w=4e-06 

m2362 1021 329 3 3 penh l=2e-06 w=1e-05 

m2363 3 1026 1025 3 penh l=2e-06 w=1.6e-05 

m2364 3 1025 1026 3 penh l=8e-06 w=4e-06 

m2365 1026 329 3 3 penh l=2e-06 w=1e-05 

m2366 1025 1026 0 0 nenh l=2e-06 w=6e-06 

m2367 0 329 1023 0 nenh l=2e-06 w=1.4e-05 

m2368 1023 697 1027 0 nenh l=2e-06 w=1e-05 

m2369 1027 151 1021 0 nenh l=2e-06 w=8e-06 

m2370 1021 699 1028 0 nenh l=2e-06 w=6e-06 

m2371 1028 146 1027 0 nenh l=2e-06 w=8e-06 

m2372 1022 699 1026 0 nenh l=2e-06 w=6e-06 

m2373 1026 692 1028 0 nenh l=2e-06 w=6e-06 

m2374 1029 697 1030 0 nenh l=2e-06 w=8e-06 

m2375 1030 146 1031 0 nenh l=2e-06 w=4e-06 

m2376 1031 694 1029 0 nenh l=2e-06 w=8e-06 

m2377 1029 699 1032 0 nenh l=2e-06 w=1e-05 

m2378 0 1030 1033 0 nenh l=2e-06 w=6e-06 

m2379 3 329 1030 3 penh l=2e-06 w=1e-05 

m2380 1030 1033 3 3 penh l=8e-06 w=4e-06 

m2381 3 1030 1033 3 penh l=2e-06 w=1.6e-05 

m2382 3 1034 1014 3 penh l=2e-06 w=1.6e-05 

m2383 3 329 1034 3 penh l=2e-06 w=1e-05 

m2384 1034 1014 3 3 penh l=8e-06 w=4e-06 

m2385 1014 1034 0 0 nenh l=2e-06 w=6e-06 

m2386 0 329 1032 0 nenh l=2e-06 w=1.4e-05 

m2387 1032 692 1035 0 nenh l=2e-06 w=1.2e-05 

m2388 1035 697 1031 0 nenh l=2e-06 w=6e-06 

m2389 1031 151 1034 0 nenh l=2e-06 w=4e-06 

m2390 1034 694 1035 0 nenh l=2e-06 w=6e-06 

m2391 1036 699 1037 0 nenh l=2e-06 w=8e-06 

m2392 1037 694 1038 0 nenh l=2e-06 w=6e-06 

m2393 1038 692 1036 0 nenh l=2e-06 w=8e-06 

m2394 1036 151 1039 0 nenh l=2e-06 w=1e-05 

m2395 0 1037 1040 0 nenh l=2e-06 w=6e-06 

m2396 3 329 1037 3 penh l=2e-06 w=1e-05 

m2397 1037 1040 3 3 penh l=8e-06 w=4e-06 

m2398 3 1037 1040 3 penh l=2e-06 w=1.6e-05 

m2399 3 1042 1041 3 penh l=2e-06 w=1.6e-05 

m2400 3 329 1042 3 penh l=2e-06 w=1e-05 

m2401 1042 1041 3 3 penh l=8e-06 w=4e-06 

m2402 1041 1042 0 0 nenh l=2e-06 w=6e-06 

m2403 0 329 1039 0 nenh l=2e-06 w=1.4e-05 

m2404 1039 146 1043 0 nenh l=2e-06 w=1e-05 

m2405 1043 692 1037 0 nenh l=2e-06 w=8e-06 

m2406 1037 697 1044 0 nenh l=2e-06 w=6e-06 

m2407 1044 699 1043 0 nenh l=2e-06 w=8e-06 

m2408 1038 697 1042 0 nenh l=2e-06 w=6e-06 

m2409 1042 694 1044 0 nenh l=2e-06 w=6e-06 

m2410 1045 697 1046 0 nenh l=2e-06 w=8e-06 

m2411 1046 151 1047 0 nenh l=2e-06 w=6e-06 

m2412 1047 694 1045 0 nenh l=2e-06 w=8e-06 

m2413 1045 692 1048 0 nenh l=2e-06 w=1e-05 

m2414 0 1046 1049 0 nenh l=2e-06 w=6e-06 

m2415 1049 1046 3 3 penh l=2e-06 w=1.6e-05 

m2416 3 1049 1046 3 penh l=8e-06 w=4e-06 

m2417 1046 329 3 3 penh l=2e-06 w=1e-05 

m2418 3 1051 1050 3 penh l=2e-06 w=1.6e-05 

m2419 3 1050 1051 3 penh l=8e-06 w=4e-06 

m2420 1051 329 3 3 penh l=2e-06 w=1e-05 

m2421 1050 1051 0 0 nenh l=2e-06 w=6e-06 

m2422 0 329 1048 0 nenh l=2e-06 w=1.4e-05 

m2423 1048 699 1052 0 nenh l=2e-06 w=1e-05 

m2424 1052 694 1046 0 nenh l=2e-06 w=8e-06 

m2425 1046 146 1053 0 nenh l=2e-06 w=6e-06 

m2426 1053 697 1052 0 nenh l=2e-06 w=8e-06 

m2427 1047 146 1051 0 nenh l=2e-06 w=6e-06 

m2428 1051 151 1053 0 nenh l=2e-06 w=6e-06 

m2429 1054 327 1055 3 penh l=2e-06 w=5e-06 

m2430 1055 329 1056 3 penh l=2e-06 w=5e-06 

m2431 1056 1057 3 3 penh l=2e-06 w=5e-06 

m2432 3 1055 1057 3 penh l=2e-06 w=6e-06 

m2433 1057 857 3 3 penh l=2e-06 w=6e-06 

m2434 3 1057 299 3 penh l=2e-06 w=2.5e-05 

m2435 1054 329 1055 0 nenh l=2e-06 w=5e-06 

m2436 1055 327 1058 0 nenh l=2e-06 w=5e-06 

m2437 1058 1057 0 0 nenh l=2e-06 w=5e-06 

m2438 0 1055 1059 0 nenh l=2e-06 w=1.3e-05 

m2439 1059 857 1057 0 nenh l=2e-06 w=1.2e-05 

m2440 0 1057 299 0 nenh l=2e-06 w=1.4e-05 

m2441 1060 126 1061 0 nenh l=2e-06 w=8e-06 

m2442 1061 729 1062 0 nenh l=2e-06 w=6e-06 

m2443 1062 131 1060 0 nenh l=2e-06 w=8e-06 

m2444 1060 731 1063 0 nenh l=2e-06 w=1e-05 

m2445 0 1061 1064 0 nenh l=2e-06 w=6e-06 

m2446 1064 1061 3 3 penh l=2e-06 w=1.6e-05 

m2447 3 1064 1061 3 penh l=8e-06 w=4e-06 

m2448 1061 329 3 3 penh l=2e-06 w=1e-05 

m2449 3 1066 1065 3 penh l=2e-06 w=1.6e-05 

m2450 3 1065 1066 3 penh l=8e-06 w=4e-06 

m2451 1066 329 3 3 penh l=2e-06 w=1e-05 

m2452 1065 1066 0 0 nenh l=2e-06 w=6e-06 

m2453 0 329 1063 0 nenh l=2e-06 w=1.4e-05 

m2454 1063 734 1067 0 nenh l=2e-06 w=1e-05 

m2455 1067 131 1061 0 nenh l=2e-06 w=8e-06 

m2456 1061 736 1068 0 nenh l=2e-06 w=6e-06 

m2457 1068 126 1067 0 nenh l=2e-06 w=8e-06 

m2458 1062 736 1066 0 nenh l=2e-06 w=6e-06 

m2459 1066 729 1068 0 nenh l=2e-06 w=6e-06 

m2460 1069 734 1070 0 nenh l=2e-06 w=8e-06 

m2461 1070 126 1071 0 nenh l=2e-06 w=4e-06 

m2462 1071 731 1069 0 nenh l=2e-06 w=8e-06 

m2463 1069 736 1072 0 nenh l=2e-06 w=1e-05 

m2464 0 1070 1073 0 nenh l=2e-06 w=6e-06 

m2465 3 329 1070 3 penh l=2e-06 w=1e-05 

m2466 1070 1073 3 3 penh l=8e-06 w=4e-06 

m2467 3 1070 1073 3 penh l=2e-06 w=1.6e-05 

m2468 3 1074 1054 3 penh l=2e-06 w=1.6e-05 

m2469 3 329 1074 3 penh l=2e-06 w=1e-05 

m2470 1074 1054 3 3 penh l=8e-06 w=4e-06 

m2471 1054 1074 0 0 nenh l=2e-06 w=6e-06 

m2472 0 329 1072 0 nenh l=2e-06 w=1.4e-05 

m2473 1072 729 1075 0 nenh l=2e-06 w=1.2e-05 

m2474 1075 734 1071 0 nenh l=2e-06 w=6e-06 

m2475 1071 131 1074 0 nenh l=2e-06 w=4e-06 

m2476 1074 731 1075 0 nenh l=2e-06 w=6e-06 

m2477 1076 736 1077 0 nenh l=2e-06 w=8e-06 

m2478 1077 731 1078 0 nenh l=2e-06 w=6e-06 

m2479 1078 729 1076 0 nenh l=2e-06 w=8e-06 

m2480 1076 131 1079 0 nenh l=2e-06 w=1e-05 

m2481 0 1077 1080 0 nenh l=2e-06 w=6e-06 

m2482 3 329 1077 3 penh l=2e-06 w=1e-05 

m2483 1077 1080 3 3 penh l=8e-06 w=4e-06 

m2484 3 1077 1080 3 penh l=2e-06 w=1.6e-05 

m2485 3 1082 1081 3 penh l=2e-06 w=1.6e-05 

m2486 3 329 1082 3 penh l=2e-06 w=1e-05 

m2487 1082 1081 3 3 penh l=8e-06 w=4e-06 

m2488 1081 1082 0 0 nenh l=2e-06 w=6e-06 

m2489 0 329 1079 0 nenh l=2e-06 w=1.4e-05 

m2490 1079 126 1083 0 nenh l=2e-06 w=1e-05 

m2491 1083 729 1077 0 nenh l=2e-06 w=8e-06 

m2492 1077 734 1084 0 nenh l=2e-06 w=6e-06 

m2493 1084 736 1083 0 nenh l=2e-06 w=8e-06 

m2494 1078 734 1082 0 nenh l=2e-06 w=6e-06 

m2495 1082 731 1084 0 nenh l=2e-06 w=6e-06 

m2496 1085 734 1086 0 nenh l=2e-06 w=8e-06 

m2497 1086 131 1087 0 nenh l=2e-06 w=6e-06 

m2498 1087 731 1085 0 nenh l=2e-06 w=8e-06 

m2499 1085 729 1088 0 nenh l=2e-06 w=1e-05 

m2500 0 1086 1089 0 nenh l=2e-06 w=6e-06 

m2501 1089 1086 3 3 penh l=2e-06 w=1.6e-05 

m2502 3 1089 1086 3 penh l=8e-06 w=4e-06 

m2503 1086 329 3 3 penh l=2e-06 w=1e-05 

m2504 3 1091 1090 3 penh l=2e-06 w=1.6e-05 

m2505 3 1090 1091 3 penh l=8e-06 w=4e-06 

m2506 1091 329 3 3 penh l=2e-06 w=1e-05 

m2507 1090 1091 0 0 nenh l=2e-06 w=6e-06 

m2508 0 329 1088 0 nenh l=2e-06 w=1.4e-05 

m2509 1088 736 1092 0 nenh l=2e-06 w=1e-05 

m2510 1092 731 1086 0 nenh l=2e-06 w=8e-06 

m2511 1086 126 1093 0 nenh l=2e-06 w=6e-06 

m2512 1093 734 1092 0 nenh l=2e-06 w=8e-06 

m2513 1087 126 1091 0 nenh l=2e-06 w=6e-06 

m2514 1091 131 1093 0 nenh l=2e-06 w=6e-06 

m2515 1094 327 1095 3 penh l=2e-06 w=5e-06 

m2516 1095 329 1096 3 penh l=2e-06 w=5e-06 

m2517 1096 1097 3 3 penh l=2e-06 w=5e-06 

m2518 3 1095 1097 3 penh l=2e-06 w=6e-06 

m2519 1097 857 3 3 penh l=2e-06 w=6e-06 

m2520 3 1097 303 3 penh l=2e-06 w=2.5e-05 

m2521 1094 329 1095 0 nenh l=2e-06 w=5e-06 

m2522 1095 327 1098 0 nenh l=2e-06 w=5e-06 

m2523 1098 1097 0 0 nenh l=2e-06 w=5e-06 

m2524 0 1095 1099 0 nenh l=2e-06 w=1.3e-05 

m2525 1099 857 1097 0 nenh l=2e-06 w=1.2e-05 

m2526 0 1097 303 0 nenh l=2e-06 w=1.4e-05 

m2527 1100 106 1101 0 nenh l=2e-06 w=8e-06 

m2528 1101 766 1102 0 nenh l=2e-06 w=6e-06 

m2529 1102 111 1100 0 nenh l=2e-06 w=8e-06 

m2530 1100 768 1103 0 nenh l=2e-06 w=1e-05 

m2531 0 1101 1104 0 nenh l=2e-06 w=6e-06 

m2532 1104 1101 3 3 penh l=2e-06 w=1.6e-05 

m2533 3 1104 1101 3 penh l=8e-06 w=4e-06 

m2534 1101 329 3 3 penh l=2e-06 w=1e-05 

m2535 3 1106 1105 3 penh l=2e-06 w=1.6e-05 

m2536 3 1105 1106 3 penh l=8e-06 w=4e-06 

m2537 1106 329 3 3 penh l=2e-06 w=1e-05 

m2538 1105 1106 0 0 nenh l=2e-06 w=6e-06 

m2539 0 329 1103 0 nenh l=2e-06 w=1.4e-05 

m2540 1103 771 1107 0 nenh l=2e-06 w=1e-05 

m2541 1107 111 1101 0 nenh l=2e-06 w=8e-06 

m2542 1101 773 1108 0 nenh l=2e-06 w=6e-06 

m2543 1108 106 1107 0 nenh l=2e-06 w=8e-06 

m2544 1102 773 1106 0 nenh l=2e-06 w=6e-06 

m2545 1106 766 1108 0 nenh l=2e-06 w=6e-06 

m2546 1109 771 1110 0 nenh l=2e-06 w=8e-06 

m2547 1110 106 1111 0 nenh l=2e-06 w=4e-06 

m2548 1111 768 1109 0 nenh l=2e-06 w=8e-06 

m2549 1109 773 1112 0 nenh l=2e-06 w=1e-05 

m2550 0 1110 1113 0 nenh l=2e-06 w=6e-06 

m2551 3 329 1110 3 penh l=2e-06 w=1e-05 

m2552 1110 1113 3 3 penh l=8e-06 w=4e-06 

m2553 3 1110 1113 3 penh l=2e-06 w=1.6e-05 

m2554 3 1114 1094 3 penh l=2e-06 w=1.6e-05 

m2555 3 329 1114 3 penh l=2e-06 w=1e-05 

m2556 1114 1094 3 3 penh l=8e-06 w=4e-06 

m2557 1094 1114 0 0 nenh l=2e-06 w=6e-06 

m2558 0 329 1112 0 nenh l=2e-06 w=1.4e-05 

m2559 1112 766 1115 0 nenh l=2e-06 w=1.2e-05 

m2560 1115 771 1111 0 nenh l=2e-06 w=6e-06 

m2561 1111 111 1114 0 nenh l=2e-06 w=4e-06 

m2562 1114 768 1115 0 nenh l=2e-06 w=6e-06 

m2563 1116 773 1117 0 nenh l=2e-06 w=8e-06 

m2564 1117 768 1118 0 nenh l=2e-06 w=6e-06 

m2565 1118 766 1116 0 nenh l=2e-06 w=8e-06 

m2566 1116 111 1119 0 nenh l=2e-06 w=1e-05 

m2567 0 1117 1120 0 nenh l=2e-06 w=6e-06 

m2568 3 329 1117 3 penh l=2e-06 w=1e-05 

m2569 1117 1120 3 3 penh l=8e-06 w=4e-06 

m2570 3 1117 1120 3 penh l=2e-06 w=1.6e-05 

m2571 3 1122 1121 3 penh l=2e-06 w=1.6e-05 

m2572 3 329 1122 3 penh l=2e-06 w=1e-05 

m2573 1122 1121 3 3 penh l=8e-06 w=4e-06 

m2574 1121 1122 0 0 nenh l=2e-06 w=6e-06 

m2575 0 329 1119 0 nenh l=2e-06 w=1.4e-05 

m2576 1119 106 1123 0 nenh l=2e-06 w=1e-05 

m2577 1123 766 1117 0 nenh l=2e-06 w=8e-06 

m2578 1117 771 1124 0 nenh l=2e-06 w=6e-06 

m2579 1124 773 1123 0 nenh l=2e-06 w=8e-06 

m2580 1118 771 1122 0 nenh l=2e-06 w=6e-06 

m2581 1122 768 1124 0 nenh l=2e-06 w=6e-06 

m2582 1125 771 1126 0 nenh l=2e-06 w=8e-06 

m2583 1126 111 1127 0 nenh l=2e-06 w=6e-06 

m2584 1127 768 1125 0 nenh l=2e-06 w=8e-06 

m2585 1125 766 1128 0 nenh l=2e-06 w=1e-05 

m2586 0 1126 1129 0 nenh l=2e-06 w=6e-06 

m2587 1129 1126 3 3 penh l=2e-06 w=1.6e-05 

m2588 3 1129 1126 3 penh l=8e-06 w=4e-06 

m2589 1126 329 3 3 penh l=2e-06 w=1e-05 

m2590 3 1131 1130 3 penh l=2e-06 w=1.6e-05 

m2591 3 1130 1131 3 penh l=8e-06 w=4e-06 

m2592 1131 329 3 3 penh l=2e-06 w=1e-05 

m2593 1130 1131 0 0 nenh l=2e-06 w=6e-06 

m2594 0 329 1128 0 nenh l=2e-06 w=1.4e-05 

m2595 1128 773 1132 0 nenh l=2e-06 w=1e-05 

m2596 1132 768 1126 0 nenh l=2e-06 w=8e-06 

m2597 1126 106 1133 0 nenh l=2e-06 w=6e-06 

m2598 1133 771 1132 0 nenh l=2e-06 w=8e-06 

m2599 1127 106 1131 0 nenh l=2e-06 w=6e-06 

m2600 1131 111 1133 0 nenh l=2e-06 w=6e-06 

m2601 1134 327 1135 3 penh l=2e-06 w=5e-06 

m2602 1135 329 1136 3 penh l=2e-06 w=5e-06 

m2603 1136 1137 3 3 penh l=2e-06 w=5e-06 

m2604 3 1135 1137 3 penh l=2e-06 w=6e-06 

m2605 1137 857 3 3 penh l=2e-06 w=6e-06 

m2606 3 1137 307 3 penh l=2e-06 w=2.5e-05 

m2607 1134 329 1135 0 nenh l=2e-06 w=5e-06 

m2608 1135 327 1138 0 nenh l=2e-06 w=5e-06 

m2609 1138 1137 0 0 nenh l=2e-06 w=5e-06 

m2610 0 1135 1139 0 nenh l=2e-06 w=1.3e-05 

m2611 1139 857 1137 0 nenh l=2e-06 w=1.2e-05 

m2612 0 1137 307 0 nenh l=2e-06 w=1.4e-05 

m2613 1140 86 1141 0 nenh l=2e-06 w=8e-06 

m2614 1141 803 1142 0 nenh l=2e-06 w=6e-06 

m2615 1142 91 1140 0 nenh l=2e-06 w=8e-06 

m2616 1140 805 1143 0 nenh l=2e-06 w=1e-05 

m2617 0 1141 1144 0 nenh l=2e-06 w=6e-06 

m2618 1144 1141 3 3 penh l=2e-06 w=1.6e-05 

m2619 3 1144 1141 3 penh l=8e-06 w=4e-06 

m2620 1141 329 3 3 penh l=2e-06 w=1e-05 

m2621 3 1146 1145 3 penh l=2e-06 w=1.6e-05 

m2622 3 1145 1146 3 penh l=8e-06 w=4e-06 

m2623 1146 329 3 3 penh l=2e-06 w=1e-05 

m2624 1145 1146 0 0 nenh l=2e-06 w=6e-06 

m2625 0 329 1143 0 nenh l=2e-06 w=1.4e-05 

m2626 1143 808 1147 0 nenh l=2e-06 w=1e-05 

m2627 1147 91 1141 0 nenh l=2e-06 w=8e-06 

m2628 1141 810 1148 0 nenh l=2e-06 w=6e-06 

m2629 1148 86 1147 0 nenh l=2e-06 w=8e-06 

m2630 1142 810 1146 0 nenh l=2e-06 w=6e-06 

m2631 1146 803 1148 0 nenh l=2e-06 w=6e-06 

m2632 1149 808 1150 0 nenh l=2e-06 w=8e-06 

m2633 1150 86 1151 0 nenh l=2e-06 w=4e-06 

m2634 1151 805 1149 0 nenh l=2e-06 w=8e-06 

m2635 1149 810 1152 0 nenh l=2e-06 w=1e-05 

m2636 0 1150 1153 0 nenh l=2e-06 w=6e-06 

m2637 3 329 1150 3 penh l=2e-06 w=1e-05 

m2638 1150 1153 3 3 penh l=8e-06 w=4e-06 

m2639 3 1150 1153 3 penh l=2e-06 w=1.6e-05 

m2640 3 1154 1134 3 penh l=2e-06 w=1.6e-05 

m2641 3 329 1154 3 penh l=2e-06 w=1e-05 

m2642 1154 1134 3 3 penh l=8e-06 w=4e-06 

m2643 1134 1154 0 0 nenh l=2e-06 w=6e-06 

m2644 0 329 1152 0 nenh l=2e-06 w=1.4e-05 

m2645 1152 803 1155 0 nenh l=2e-06 w=1.2e-05 

m2646 1155 808 1151 0 nenh l=2e-06 w=6e-06 

m2647 1151 91 1154 0 nenh l=2e-06 w=4e-06 

m2648 1154 805 1155 0 nenh l=2e-06 w=6e-06 

m2649 1156 810 1157 0 nenh l=2e-06 w=8e-06 

m2650 1157 805 1158 0 nenh l=2e-06 w=6e-06 

m2651 1158 803 1156 0 nenh l=2e-06 w=8e-06 

m2652 1156 91 1159 0 nenh l=2e-06 w=1e-05 

m2653 0 1157 1160 0 nenh l=2e-06 w=6e-06 

m2654 3 329 1157 3 penh l=2e-06 w=1e-05 

m2655 1157 1160 3 3 penh l=8e-06 w=4e-06 

m2656 3 1157 1160 3 penh l=2e-06 w=1.6e-05 

m2657 3 1162 1161 3 penh l=2e-06 w=1.6e-05 

m2658 3 329 1162 3 penh l=2e-06 w=1e-05 

m2659 1162 1161 3 3 penh l=8e-06 w=4e-06 

m2660 1161 1162 0 0 nenh l=2e-06 w=6e-06 

m2661 0 329 1159 0 nenh l=2e-06 w=1.4e-05 

m2662 1159 86 1163 0 nenh l=2e-06 w=1e-05 

m2663 1163 803 1157 0 nenh l=2e-06 w=8e-06 

m2664 1157 808 1164 0 nenh l=2e-06 w=6e-06 

m2665 1164 810 1163 0 nenh l=2e-06 w=8e-06 

m2666 1158 808 1162 0 nenh l=2e-06 w=6e-06 

m2667 1162 805 1164 0 nenh l=2e-06 w=6e-06 

m2668 1165 808 1166 0 nenh l=2e-06 w=8e-06 

m2669 1166 91 1167 0 nenh l=2e-06 w=6e-06 

m2670 1167 805 1165 0 nenh l=2e-06 w=8e-06 

m2671 1165 803 1168 0 nenh l=2e-06 w=1e-05 

m2672 0 1166 1169 0 nenh l=2e-06 w=6e-06 

m2673 1169 1166 3 3 penh l=2e-06 w=1.6e-05 

m2674 3 1169 1166 3 penh l=8e-06 w=4e-06 

m2675 1166 329 3 3 penh l=2e-06 w=1e-05 

m2676 3 1171 1170 3 penh l=2e-06 w=1.6e-05 

m2677 3 1170 1171 3 penh l=8e-06 w=4e-06 

m2678 1171 329 3 3 penh l=2e-06 w=1e-05 

m2679 1170 1171 0 0 nenh l=2e-06 w=6e-06 

m2680 0 329 1168 0 nenh l=2e-06 w=1.4e-05 

m2681 1168 810 1172 0 nenh l=2e-06 w=1e-05 

m2682 1172 805 1166 0 nenh l=2e-06 w=8e-06 

m2683 1166 86 1173 0 nenh l=2e-06 w=6e-06 

m2684 1173 808 1172 0 nenh l=2e-06 w=8e-06 

m2685 1167 86 1171 0 nenh l=2e-06 w=6e-06 

m2686 1171 91 1173 0 nenh l=2e-06 w=6e-06 

m2687 1174 1009 1175 0 nenh l=2e-06 w=1.2e-05 

m2688 1174 969 1176 0 nenh l=2e-06 w=1.2e-05 

m2689 1176 929 1177 0 nenh l=2e-06 w=1.2e-05 

m2690 1177 889 1178 0 nenh l=2e-06 w=1.4e-05 

m2691 0 1175 1179 0 nenh l=2e-06 w=6e-06 

m2692 3 329 1175 3 penh l=2e-06 w=1e-05 

m2693 1175 1179 3 3 penh l=8e-06 w=4e-06 

m2694 3 1175 1179 3 penh l=2e-06 w=1.6e-05 

m2695 3 1181 1180 3 penh l=2e-06 w=1.6e-05 

m2696 3 329 1181 3 penh l=2e-06 w=1e-05 

m2697 1181 1180 3 3 penh l=8e-06 w=4e-06 

m2698 1180 1181 0 0 nenh l=2e-06 w=6e-06 

m2699 0 329 1178 0 nenh l=2e-06 w=1.4e-05 

m2700 1182 930 1178 0 nenh l=2e-06 w=8e-06 

m2701 1178 969 1183 0 nenh l=2e-06 w=1e-05 

m2702 1183 1010 1184 0 nenh l=2e-06 w=1e-05 

m2703 1184 970 1178 0 nenh l=2e-06 w=8e-06 

m2704 1178 890 1181 0 nenh l=2e-06 w=6e-06 

m2705 1181 889 1182 0 nenh l=2e-06 w=6e-06 

m2706 1182 929 1184 0 nenh l=2e-06 w=8e-06 

m2707 1185 1000 1186 0 nenh l=2e-06 w=1.2e-05 

m2708 1185 960 1187 0 nenh l=2e-06 w=1.2e-05 

m2709 1187 920 1188 0 nenh l=2e-06 w=1.2e-05 

m2710 1188 880 1189 0 nenh l=2e-06 w=1.4e-05 

m2711 0 1186 1190 0 nenh l=2e-06 w=6e-06 

m2712 3 329 1186 3 penh l=2e-06 w=1e-05 

m2713 1186 1190 3 3 penh l=8e-06 w=4e-06 

m2714 3 1186 1190 3 penh l=2e-06 w=1.6e-05 

m2715 3 1192 1191 3 penh l=2e-06 w=1.6e-05 

m2716 3 329 1192 3 penh l=2e-06 w=1e-05 

m2717 1192 1191 3 3 penh l=8e-06 w=4e-06 

m2718 1191 1192 0 0 nenh l=2e-06 w=6e-06 

m2719 0 329 1189 0 nenh l=2e-06 w=1.4e-05 

m2720 1193 921 1189 0 nenh l=2e-06 w=8e-06 

m2721 1189 960 1194 0 nenh l=2e-06 w=1e-05 

m2722 1194 1001 1195 0 nenh l=2e-06 w=1e-05 

m2723 1195 961 1189 0 nenh l=2e-06 w=8e-06 

m2724 1189 881 1192 0 nenh l=2e-06 w=6e-06 

m2725 1192 880 1193 0 nenh l=2e-06 w=6e-06 

m2726 1193 920 1195 0 nenh l=2e-06 w=8e-06 

m2727 1196 984 1197 0 nenh l=2e-06 w=1.2e-05 

m2728 1196 944 1198 0 nenh l=2e-06 w=1.2e-05 

m2729 1198 904 1199 0 nenh l=2e-06 w=1.2e-05 

m2730 1199 864 1200 0 nenh l=2e-06 w=1.4e-05 

m2731 0 1197 1201 0 nenh l=2e-06 w=6e-06 

m2732 3 329 1197 3 penh l=2e-06 w=1e-05 

m2733 1197 1201 3 3 penh l=8e-06 w=4e-06 

m2734 3 1197 1201 3 penh l=2e-06 w=1.6e-05 

m2735 3 1203 1202 3 penh l=2e-06 w=1.6e-05 

m2736 3 329 1203 3 penh l=2e-06 w=1e-05 

m2737 1203 1202 3 3 penh l=8e-06 w=4e-06 

m2738 1202 1203 0 0 nenh l=2e-06 w=6e-06 

m2739 0 329 1200 0 nenh l=2e-06 w=1.4e-05 

m2740 1204 905 1200 0 nenh l=2e-06 w=8e-06 

m2741 1200 944 1205 0 nenh l=2e-06 w=1e-05 

m2742 1205 985 1206 0 nenh l=2e-06 w=1e-05 

m2743 1206 945 1200 0 nenh l=2e-06 w=8e-06 

m2744 1200 865 1203 0 nenh l=2e-06 w=6e-06 

m2745 1203 864 1204 0 nenh l=2e-06 w=6e-06 

m2746 1204 904 1206 0 nenh l=2e-06 w=8e-06 

m2747 1207 953 1208 0 nenh l=2e-06 w=8e-06 

m2748 1208 913 1209 0 nenh l=2e-06 w=6e-06 

m2749 1209 274 1210 0 nenh l=2e-06 w=5e-06 

m2750 1210 873 1211 0 nenh l=2e-06 w=5e-06 

m2751 1211 280 1208 0 nenh l=2e-06 w=6e-06 

m2752 1208 285 1212 0 nenh l=2e-06 w=8e-06 

m2753 1212 993 1213 0 nenh l=2e-06 w=1e-05 

m2754 0 1210 1214 0 nenh l=2e-06 w=6e-06 

m2755 3 329 1210 3 penh l=2e-06 w=1.6e-05 

m2756 1210 1214 3 3 penh l=8e-06 w=4e-06 

m2757 3 1210 1214 3 penh l=2e-06 w=1.6e-05 

m2758 3 1216 1215 3 penh l=2e-06 w=1.6e-05 

m2759 3 329 1216 3 penh l=2e-06 w=1.6e-05 

m2760 1216 1215 3 3 penh l=8e-06 w=4e-06 

m2761 1215 1216 0 0 nenh l=2e-06 w=6e-06 

m2762 0 329 1213 0 nenh l=2e-06 w=4e-06 

m2763 1213 290 1207 0 nenh l=2e-06 w=1e-05 

m2764 1207 285 1217 0 nenh l=2e-06 w=8e-06 

m2765 1217 280 1209 0 nenh l=2e-06 w=7e-06 

m2766 1209 873 1216 0 nenh l=2e-06 w=6e-06 

m2767 1216 274 1211 0 nenh l=2e-06 w=6e-06 

m2768 1211 913 1217 0 nenh l=2e-06 w=7e-06 

m2769 1217 953 1212 0 nenh l=2e-06 w=8e-06 

m2770 1218 1073 1219 0 nenh l=2e-06 w=8e-06 

m2771 1219 1113 1220 0 nenh l=2e-06 w=6e-06 

m2772 1220 307 1221 0 nenh l=2e-06 w=5e-06 

m2773 1221 1153 1222 0 nenh l=2e-06 w=5e-06 

m2774 1222 303 1219 0 nenh l=2e-06 w=6e-06 

m2775 1219 299 1223 0 nenh l=2e-06 w=8e-06 

m2776 1223 1033 1224 0 nenh l=2e-06 w=1e-05 

m2777 0 1221 1225 0 nenh l=2e-06 w=6e-06 

m2778 3 329 1221 3 penh l=2e-06 w=1.6e-05 

m2779 1221 1225 3 3 penh l=8e-06 w=4e-06 

m2780 3 1221 1225 3 penh l=2e-06 w=1.6e-05 

m2781 3 1227 1226 3 penh l=2e-06 w=1.6e-05 

m2782 3 329 1227 3 penh l=2e-06 w=1.6e-05 

m2783 1227 1226 3 3 penh l=8e-06 w=4e-06 

m2784 1226 1227 0 0 nenh l=2e-06 w=6e-06 

m2785 0 329 1224 0 nenh l=2e-06 w=4e-06 

m2786 1224 295 1218 0 nenh l=2e-06 w=1e-05 

m2787 1218 299 1228 0 nenh l=2e-06 w=8e-06 

m2788 1228 303 1220 0 nenh l=2e-06 w=7e-06 

m2789 1220 1153 1227 0 nenh l=2e-06 w=6e-06 

m2790 1227 307 1222 0 nenh l=2e-06 w=6e-06 

m2791 1222 1113 1228 0 nenh l=2e-06 w=7e-06 

m2792 1228 1073 1223 0 nenh l=2e-06 w=8e-06 

m2793 1229 1179 1230 0 nenh l=2e-06 w=6e-06 

m2794 1230 1232 1231 0 nenh l=2e-06 w=6e-06 

m2795 0 1229 1233 0 nenh l=2e-06 w=6e-06 

m2796 3 329 1229 3 penh l=2e-06 w=1e-05 

m2797 1229 1233 3 3 penh l=8e-06 w=4e-06 

m2798 3 1229 1233 3 penh l=2e-06 w=1.6e-05 

m2799 3 1235 1234 3 penh l=2e-06 w=1.6e-05 

m2800 3 329 1235 3 penh l=2e-06 w=1e-05 

m2801 1235 1234 3 3 penh l=8e-06 w=4e-06 

m2802 1234 1235 0 0 nenh l=2e-06 w=6e-06 

m2803 0 329 1231 0 nenh l=2e-06 w=1.2e-05 

m2804 1231 1237 1236 0 nenh l=2e-06 w=6e-06 

m2805 1236 1179 1235 0 nenh l=2e-06 w=6e-06 

m2806 1235 1180 1231 0 nenh l=2e-06 w=6e-06 

m2807 1238 1190 1239 0 nenh l=2e-06 w=6e-06 

m2808 1239 1241 1240 0 nenh l=2e-06 w=6e-06 

m2809 0 1238 1242 0 nenh l=2e-06 w=6e-06 

m2810 3 329 1238 3 penh l=2e-06 w=1e-05 

m2811 1238 1242 3 3 penh l=8e-06 w=4e-06 

m2812 3 1238 1242 3 penh l=2e-06 w=1.6e-05 

m2813 3 1244 1243 3 penh l=2e-06 w=1.6e-05 

m2814 3 329 1244 3 penh l=2e-06 w=1e-05 

m2815 1244 1243 3 3 penh l=8e-06 w=4e-06 

m2816 1243 1244 0 0 nenh l=2e-06 w=6e-06 

m2817 0 329 1240 0 nenh l=2e-06 w=1.2e-05 

m2818 1240 1246 1245 0 nenh l=2e-06 w=6e-06 

m2819 1245 1190 1244 0 nenh l=2e-06 w=6e-06 

m2820 1244 1191 1240 0 nenh l=2e-06 w=6e-06 

m2821 1247 1201 1248 0 nenh l=2e-06 w=6e-06 

m2822 1248 1250 1249 0 nenh l=2e-06 w=6e-06 

m2823 0 1247 1251 0 nenh l=2e-06 w=6e-06 

m2824 3 329 1247 3 penh l=2e-06 w=1e-05 

m2825 1247 1251 3 3 penh l=8e-06 w=4e-06 

m2826 3 1247 1251 3 penh l=2e-06 w=1.6e-05 

m2827 3 1253 1252 3 penh l=2e-06 w=1.6e-05 

m2828 3 329 1253 3 penh l=2e-06 w=1e-05 

m2829 1253 1252 3 3 penh l=8e-06 w=4e-06 

m2830 1252 1253 0 0 nenh l=2e-06 w=6e-06 

m2831 0 329 1249 0 nenh l=2e-06 w=1.2e-05 

m2832 1249 1255 1254 0 nenh l=2e-06 w=6e-06 

m2833 1254 1201 1253 0 nenh l=2e-06 w=6e-06 

m2834 1253 1202 1249 0 nenh l=2e-06 w=6e-06 

m2835 1256 1215 1257 0 nenh l=2e-06 w=4e-06 

m2836 1257 1214 1258 0 nenh l=2e-06 w=4e-06 

m2837 0 1257 1259 0 nenh l=2e-06 w=6e-06 

m2838 3 329 1257 3 penh l=2e-06 w=1.6e-05 

m2839 1257 1259 3 3 penh l=8e-06 w=4e-06 

m2840 3 1257 1259 3 penh l=2e-06 w=1.6e-05 

m2841 3 1261 1260 3 penh l=2e-06 w=1.6e-05 

m2842 3 329 1261 3 penh l=2e-06 w=1.6e-05 

m2843 1261 1260 3 3 penh l=8e-06 w=4e-06 

m2844 1260 1261 0 0 nenh l=2e-06 w=6e-06 

m2845 0 329 1262 0 nenh l=2e-06 w=4e-06 

m2846 1262 1226 1256 0 nenh l=2e-06 w=8e-06 

m2847 1256 1214 1261 0 nenh l=2e-06 w=4e-06 

m2848 1261 1215 1258 0 nenh l=2e-06 w=4e-06 

m2849 1258 1225 1262 0 nenh l=2e-06 w=8e-06 

m2850 1263 1242 1264 0 nenh l=2e-06 w=8e-06 

m2851 1264 1259 1265 0 nenh l=2e-06 w=6e-06 

m2852 1265 1234 1266 0 nenh l=2e-06 w=5e-06 

m2853 1266 1233 1267 0 nenh l=2e-06 w=5e-06 

m2854 1267 1260 1264 0 nenh l=2e-06 w=6e-06 

m2855 1264 1243 1268 0 nenh l=2e-06 w=8e-06 

m2856 1268 1251 1269 0 nenh l=2e-06 w=1e-05 

m2857 0 1266 1270 0 nenh l=2e-06 w=6e-06 

m2858 3 329 1266 3 penh l=2e-06 w=1.6e-05 

m2859 1266 1270 3 3 penh l=8e-06 w=4e-06 

m2860 3 1266 1270 3 penh l=2e-06 w=1.6e-05 

m2861 3 1272 1271 3 penh l=2e-06 w=1.6e-05 

m2862 3 329 1272 3 penh l=2e-06 w=1.6e-05 

m2863 1272 1271 3 3 penh l=8e-06 w=4e-06 

m2864 1271 1272 0 0 nenh l=2e-06 w=6e-06 

m2865 0 329 1269 0 nenh l=2e-06 w=4e-06 

m2866 1269 1252 1263 0 nenh l=2e-06 w=1e-05 

m2867 1263 1243 1273 0 nenh l=2e-06 w=8e-06 

m2868 1273 1260 1265 0 nenh l=2e-06 w=7e-06 

m2869 1265 1233 1272 0 nenh l=2e-06 w=6e-06 

m2870 1272 1234 1267 0 nenh l=2e-06 w=6e-06 

m2871 1267 1259 1273 0 nenh l=2e-06 w=7e-06 

m2872 1273 1242 1268 0 nenh l=2e-06 w=8e-06 

m2873 1274 1169 1275 0 nenh l=2e-06 w=1.2e-05 

m2874 1274 1129 1276 0 nenh l=2e-06 w=1.2e-05 

m2875 1276 1049 1277 0 nenh l=2e-06 w=1.2e-05 

m2876 1277 1089 1278 0 nenh l=2e-06 w=1.4e-05 

m2877 0 1275 1232 0 nenh l=2e-06 w=6e-06 

m2878 3 329 1275 3 penh l=2e-06 w=1e-05 

m2879 1275 1232 3 3 penh l=8e-06 w=4e-06 

m2880 3 1275 1232 3 penh l=2e-06 w=1.6e-05 

m2881 3 1279 1237 3 penh l=2e-06 w=1.6e-05 

m2882 3 329 1279 3 penh l=2e-06 w=1e-05 

m2883 1279 1237 3 3 penh l=8e-06 w=4e-06 

m2884 1237 1279 0 0 nenh l=2e-06 w=6e-06 

m2885 0 329 1278 0 nenh l=2e-06 w=1.4e-05 

m2886 1280 1050 1278 0 nenh l=2e-06 w=8e-06 

m2887 1278 1129 1281 0 nenh l=2e-06 w=1e-05 

m2888 1281 1170 1282 0 nenh l=2e-06 w=1e-05 

m2889 1282 1130 1278 0 nenh l=2e-06 w=8e-06 

m2890 1278 1090 1279 0 nenh l=2e-06 w=6e-06 

m2891 1279 1089 1280 0 nenh l=2e-06 w=6e-06 

m2892 1280 1049 1282 0 nenh l=2e-06 w=8e-06 

m2893 1283 1040 1284 0 nenh l=2e-06 w=1.2e-05 

m2894 1283 1080 1285 0 nenh l=2e-06 w=1.2e-05 

m2895 1285 1120 1286 0 nenh l=2e-06 w=1.2e-05 

m2896 1286 1160 1287 0 nenh l=2e-06 w=1.4e-05 

m2897 0 1284 1241 0 nenh l=2e-06 w=6e-06 

m2898 3 329 1284 3 penh l=2e-06 w=1e-05 

m2899 1284 1241 3 3 penh l=8e-06 w=4e-06 

m2900 3 1284 1241 3 penh l=2e-06 w=1.6e-05 

m2901 3 1288 1246 3 penh l=2e-06 w=1.6e-05 

m2902 3 329 1288 3 penh l=2e-06 w=1e-05 

m2903 1288 1246 3 3 penh l=8e-06 w=4e-06 

m2904 1246 1288 0 0 nenh l=2e-06 w=6e-06 

m2905 0 329 1287 0 nenh l=2e-06 w=1.4e-05 

m2906 1289 1121 1287 0 nenh l=2e-06 w=8e-06 

m2907 1287 1080 1290 0 nenh l=2e-06 w=1e-05 

m2908 1290 1041 1291 0 nenh l=2e-06 w=1e-05 

m2909 1291 1081 1287 0 nenh l=2e-06 w=8e-06 

m2910 1287 1161 1288 0 nenh l=2e-06 w=6e-06 

m2911 1288 1160 1289 0 nenh l=2e-06 w=6e-06 

m2912 1289 1120 1291 0 nenh l=2e-06 w=8e-06 

m2913 1292 1024 1293 0 nenh l=2e-06 w=1.2e-05 

m2914 1292 1064 1294 0 nenh l=2e-06 w=1.2e-05 

m2915 1294 1104 1295 0 nenh l=2e-06 w=1.2e-05 

m2916 1295 1144 1296 0 nenh l=2e-06 w=1.4e-05 

m2917 0 1293 1250 0 nenh l=2e-06 w=6e-06 

m2918 3 329 1293 3 penh l=2e-06 w=1e-05 

m2919 1293 1250 3 3 penh l=8e-06 w=4e-06 

m2920 3 1293 1250 3 penh l=2e-06 w=1.6e-05 

m2921 3 1297 1255 3 penh l=2e-06 w=1.6e-05 

m2922 3 329 1297 3 penh l=2e-06 w=1e-05 

m2923 1297 1255 3 3 penh l=8e-06 w=4e-06 

m2924 1255 1297 0 0 nenh l=2e-06 w=6e-06 

m2925 0 329 1296 0 nenh l=2e-06 w=1.4e-05 

m2926 1298 1105 1296 0 nenh l=2e-06 w=8e-06 

m2927 1296 1064 1299 0 nenh l=2e-06 w=1e-05 

m2928 1299 1025 1300 0 nenh l=2e-06 w=1e-05 

m2929 1300 1065 1296 0 nenh l=2e-06 w=8e-06 

m2930 1296 1145 1297 0 nenh l=2e-06 w=6e-06 

m2931 1297 1144 1298 0 nenh l=2e-06 w=6e-06 

m2932 1298 1104 1300 0 nenh l=2e-06 w=8e-06 

m2933 1234 327 1301 3 penh l=2e-06 w=5e-06 

m2934 1301 329 1302 3 penh l=2e-06 w=5e-06 

m2935 1302 1303 3 3 penh l=2e-06 w=5e-06 

m2936 3 1301 1303 3 penh l=2e-06 w=6e-06 

m2937 1303 857 3 3 penh l=2e-06 w=6e-06 

m2938 3 1303 311 3 penh l=2e-06 w=2.5e-05 

m2939 1234 329 1301 0 nenh l=2e-06 w=5e-06 

m2940 1301 327 1304 0 nenh l=2e-06 w=5e-06 

m2941 1304 1303 0 0 nenh l=2e-06 w=5e-06 

m2942 0 1301 1305 0 nenh l=2e-06 w=1.3e-05 

m2943 1305 857 1303 0 nenh l=2e-06 w=1.2e-05 

m2944 0 1303 311 0 nenh l=2e-06 w=1.4e-05 

m2945 1243 327 1306 3 penh l=2e-06 w=5e-06 

m2946 1306 329 1307 3 penh l=2e-06 w=5e-06 

m2947 1307 1308 3 3 penh l=2e-06 w=5e-06 

m2948 3 1306 1308 3 penh l=2e-06 w=6e-06 

m2949 1308 857 3 3 penh l=2e-06 w=6e-06 

m2950 3 1308 315 3 penh l=2e-06 w=2.5e-05 

m2951 1243 329 1306 0 nenh l=2e-06 w=5e-06 

m2952 1306 327 1309 0 nenh l=2e-06 w=5e-06 

m2953 1309 1308 0 0 nenh l=2e-06 w=5e-06 

m2954 0 1306 1310 0 nenh l=2e-06 w=1.3e-05 

m2955 1310 857 1308 0 nenh l=2e-06 w=1.2e-05 

m2956 0 1308 315 0 nenh l=2e-06 w=1.4e-05 

m2957 1252 327 1311 3 penh l=2e-06 w=5e-06 

m2958 1311 329 1312 3 penh l=2e-06 w=5e-06 

m2959 1312 1313 3 3 penh l=2e-06 w=5e-06 

m2960 3 1311 1313 3 penh l=2e-06 w=6e-06 

m2961 1313 857 3 3 penh l=2e-06 w=6e-06 

m2962 3 1313 319 3 penh l=2e-06 w=2.5e-05 

m2963 1252 329 1311 0 nenh l=2e-06 w=5e-06 

m2964 1311 327 1314 0 nenh l=2e-06 w=5e-06 

m2965 1314 1313 0 0 nenh l=2e-06 w=5e-06 

m2966 0 1311 1315 0 nenh l=2e-06 w=1.3e-05 

m2967 1315 857 1313 0 nenh l=2e-06 w=1.2e-05 

m2968 0 1313 319 0 nenh l=2e-06 w=1.4e-05 

m2969 1271 327 1316 3 penh l=2e-06 w=5e-06 

m2970 1316 329 1317 3 penh l=2e-06 w=5e-06 

m2971 1317 1318 3 3 penh l=2e-06 w=5e-06 

m2972 3 1316 1318 3 penh l=2e-06 w=6e-06 

m2973 1318 857 3 3 penh l=2e-06 w=6e-06 

m2974 3 1318 1319 3 penh l=2e-06 w=2.5e-05 

m2975 1271 329 1316 0 nenh l=2e-06 w=5e-06 

m2976 1316 327 1320 0 nenh l=2e-06 w=5e-06 

m2977 1320 1318 0 0 nenh l=2e-06 w=5e-06 

m2978 0 1316 1321 0 nenh l=2e-06 w=1.3e-05 

m2979 1321 857 1318 0 nenh l=2e-06 w=1.2e-05 

m2980 0 1318 1319 0 nenh l=2e-06 w=1.4e-05 

m2981 1270 327 1322 3 penh l=2e-06 w=5e-06 

m2982 1322 329 1323 3 penh l=2e-06 w=5e-06 

m2983 1323 1324 3 3 penh l=2e-06 w=5e-06 

m2984 3 1322 1324 3 penh l=2e-06 w=6e-06 

m2985 1324 857 3 3 penh l=2e-06 w=6e-06 

m2986 3 1324 1325 3 penh l=2e-06 w=2.5e-05 

m2987 1270 329 1322 0 nenh l=2e-06 w=5e-06 

m2988 1322 327 1326 0 nenh l=2e-06 w=5e-06 

m2989 1326 1324 0 0 nenh l=2e-06 w=5e-06 

m2990 0 1322 1327 0 nenh l=2e-06 w=1.3e-05 

m2991 1327 857 1324 0 nenh l=2e-06 w=1.2e-05 

m2992 0 1324 1325 0 nenh l=2e-06 w=1.4e-05 

m2993 75 1329 1328 3 penh l=2e-06 w=6e-06 

m2994 1328 1331 1330 3 penh l=2e-06 w=6e-06 

m2995 1328 81 1332 3 penh l=2e-06 w=6e-06 

m2996 1332 83 1333 3 penh l=2e-06 w=6e-06 

m2997 1333 1334 3 3 penh l=2e-06 w=6e-06 

m2998 3 1332 1334 3 penh l=2e-06 w=6e-06 

m2999 1334 74 3 3 penh l=2e-06 w=6e-06 

m3000 3 1334 1330 3 penh l=2e-06 w=6e-06 

m3001 3 1330 1335 3 penh l=2e-06 w=2.4e-05 

m3002 75 1331 1328 0 nenh l=2e-06 w=4e-06 

m3003 1328 1329 1330 0 nenh l=2e-06 w=4e-06 

m3004 3 1335 808 3 penh l=2e-06 w=2.8e-05 

m3005 808 1335 3 3 penh l=2e-06 w=3e-05 

m3006 808 1335 3 3 penh l=2e-06 w=1.8e-05 

m3007 1328 83 1332 0 nenh l=2e-06 w=4e-06 

m3008 1332 81 1336 0 nenh l=2e-06 w=4e-06 

m3009 1336 1334 0 0 nenh l=2e-06 w=4e-06 

m3010 0 1332 1337 0 nenh l=2e-06 w=8e-06 

m3011 1337 74 1334 0 nenh l=2e-06 w=8e-06 

m3012 3 1335 808 3 penh l=2e-06 w=1.8e-05 

m3013 1330 1334 0 0 nenh l=2e-06 w=4e-06 

m3014 0 1330 1335 0 nenh l=2e-06 w=1.6e-05 

m3015 808 1335 0 0 nenh l=2e-06 w=1.4e-05 

m3016 0 1335 808 0 nenh l=2e-06 w=3.1e-05 

m3017 808 1335 0 0 nenh l=2e-06 w=1.9e-05 

m3018 0 1339 1338 0 nenh l=2e-06 w=1.6e-05 

m3019 0 1338 805 0 nenh l=2e-06 w=3.1e-05 

m3020 92 1331 1340 0 nenh l=2e-06 w=4e-06 

m3021 1340 1329 1339 0 nenh l=2e-06 w=4e-06 

m3022 1340 83 1341 0 nenh l=2e-06 w=4e-06 

m3023 1341 81 1342 0 nenh l=2e-06 w=4e-06 

m3024 1342 1343 0 0 nenh l=2e-06 w=4e-06 

m3025 0 1341 1344 0 nenh l=2e-06 w=8e-06 

m3026 1344 74 1343 0 nenh l=2e-06 w=8e-06 

m3027 1339 1343 0 0 nenh l=2e-06 w=4e-06 

m3028 0 1338 805 0 nenh l=2e-06 w=1.4e-05 

m3029 805 1338 0 0 nenh l=2e-06 w=1.9e-05 

m3030 92 1329 1340 3 penh l=2e-06 w=6e-06 

m3031 1340 1331 1339 3 penh l=2e-06 w=6e-06 

m3032 1340 81 1341 3 penh l=2e-06 w=6e-06 

m3033 1341 83 1345 3 penh l=2e-06 w=6e-06 

m3034 1345 1343 3 3 penh l=2e-06 w=6e-06 

m3035 3 1341 1343 3 penh l=2e-06 w=6e-06 

m3036 1343 74 3 3 penh l=2e-06 w=6e-06 

m3037 3 1343 1339 3 penh l=2e-06 w=6e-06 

m3038 3 1339 1338 3 penh l=2e-06 w=2.4e-05 

m3039 3 1338 805 3 penh l=2e-06 w=1.8e-05 

m3040 805 1338 3 3 penh l=2e-06 w=3e-05 

m3041 3 1338 805 3 penh l=2e-06 w=1.8e-05 

m3042 805 1338 3 3 penh l=2e-06 w=2.8e-05 

m3043 99 1329 1346 3 penh l=2e-06 w=6e-06 

m3044 1346 1331 1347 3 penh l=2e-06 w=6e-06 

m3045 1346 81 1348 3 penh l=2e-06 w=6e-06 

m3046 1348 83 1349 3 penh l=2e-06 w=6e-06 

m3047 1349 1350 3 3 penh l=2e-06 w=6e-06 

m3048 3 1348 1350 3 penh l=2e-06 w=6e-06 

m3049 1350 74 3 3 penh l=2e-06 w=6e-06 

m3050 3 1350 1347 3 penh l=2e-06 w=6e-06 

m3051 3 1347 1351 3 penh l=2e-06 w=2.4e-05 

m3052 99 1331 1346 0 nenh l=2e-06 w=4e-06 

m3053 1346 1329 1347 0 nenh l=2e-06 w=4e-06 

m3054 3 1351 771 3 penh l=2e-06 w=2.8e-05 

m3055 771 1351 3 3 penh l=2e-06 w=3e-05 

m3056 771 1351 3 3 penh l=2e-06 w=1.8e-05 

m3057 1346 83 1348 0 nenh l=2e-06 w=4e-06 

m3058 1348 81 1352 0 nenh l=2e-06 w=4e-06 

m3059 1352 1350 0 0 nenh l=2e-06 w=4e-06 

m3060 0 1348 1353 0 nenh l=2e-06 w=8e-06 

m3061 1353 74 1350 0 nenh l=2e-06 w=8e-06 

m3062 3 1351 771 3 penh l=2e-06 w=1.8e-05 

m3063 1347 1350 0 0 nenh l=2e-06 w=4e-06 

m3064 0 1347 1351 0 nenh l=2e-06 w=1.6e-05 

m3065 771 1351 0 0 nenh l=2e-06 w=1.4e-05 

m3066 0 1351 771 0 nenh l=2e-06 w=3.1e-05 

m3067 771 1351 0 0 nenh l=2e-06 w=1.9e-05 

m3068 0 1355 1354 0 nenh l=2e-06 w=1.6e-05 

m3069 0 1354 768 0 nenh l=2e-06 w=3.1e-05 

m3070 112 1331 1356 0 nenh l=2e-06 w=4e-06 

m3071 1356 1329 1355 0 nenh l=2e-06 w=4e-06 

m3072 1356 83 1357 0 nenh l=2e-06 w=4e-06 

m3073 1357 81 1358 0 nenh l=2e-06 w=4e-06 

m3074 1358 1359 0 0 nenh l=2e-06 w=4e-06 

m3075 0 1357 1360 0 nenh l=2e-06 w=8e-06 

m3076 1360 74 1359 0 nenh l=2e-06 w=8e-06 

m3077 1355 1359 0 0 nenh l=2e-06 w=4e-06 

m3078 0 1354 768 0 nenh l=2e-06 w=1.4e-05 

m3079 768 1354 0 0 nenh l=2e-06 w=1.9e-05 

m3080 112 1329 1356 3 penh l=2e-06 w=6e-06 

m3081 1356 1331 1355 3 penh l=2e-06 w=6e-06 

m3082 1356 81 1357 3 penh l=2e-06 w=6e-06 

m3083 1357 83 1361 3 penh l=2e-06 w=6e-06 

m3084 1361 1359 3 3 penh l=2e-06 w=6e-06 

m3085 3 1357 1359 3 penh l=2e-06 w=6e-06 

m3086 1359 74 3 3 penh l=2e-06 w=6e-06 

m3087 3 1359 1355 3 penh l=2e-06 w=6e-06 

m3088 3 1355 1354 3 penh l=2e-06 w=2.4e-05 

m3089 3 1354 768 3 penh l=2e-06 w=1.8e-05 

m3090 768 1354 3 3 penh l=2e-06 w=3e-05 

m3091 3 1354 768 3 penh l=2e-06 w=1.8e-05 

m3092 768 1354 3 3 penh l=2e-06 w=2.8e-05 

m3093 119 1329 1362 3 penh l=2e-06 w=6e-06 

m3094 1362 1331 1363 3 penh l=2e-06 w=6e-06 

m3095 1362 81 1364 3 penh l=2e-06 w=6e-06 

m3096 1364 83 1365 3 penh l=2e-06 w=6e-06 

m3097 1365 1366 3 3 penh l=2e-06 w=6e-06 

m3098 3 1364 1366 3 penh l=2e-06 w=6e-06 

m3099 1366 74 3 3 penh l=2e-06 w=6e-06 

m3100 3 1366 1363 3 penh l=2e-06 w=6e-06 

m3101 3 1363 1367 3 penh l=2e-06 w=2.4e-05 

m3102 119 1331 1362 0 nenh l=2e-06 w=4e-06 

m3103 1362 1329 1363 0 nenh l=2e-06 w=4e-06 

m3104 3 1367 734 3 penh l=2e-06 w=2.8e-05 

m3105 734 1367 3 3 penh l=2e-06 w=3e-05 

m3106 734 1367 3 3 penh l=2e-06 w=1.8e-05 

m3107 1362 83 1364 0 nenh l=2e-06 w=4e-06 

m3108 1364 81 1368 0 nenh l=2e-06 w=4e-06 

m3109 1368 1366 0 0 nenh l=2e-06 w=4e-06 

m3110 0 1364 1369 0 nenh l=2e-06 w=8e-06 

m3111 1369 74 1366 0 nenh l=2e-06 w=8e-06 

m3112 3 1367 734 3 penh l=2e-06 w=1.8e-05 

m3113 1363 1366 0 0 nenh l=2e-06 w=4e-06 

m3114 0 1363 1367 0 nenh l=2e-06 w=1.6e-05 

m3115 734 1367 0 0 nenh l=2e-06 w=1.4e-05 

m3116 0 1367 734 0 nenh l=2e-06 w=3.1e-05 

m3117 734 1367 0 0 nenh l=2e-06 w=1.9e-05 

m3118 0 1371 1370 0 nenh l=2e-06 w=1.6e-05 

m3119 0 1370 731 0 nenh l=2e-06 w=3.1e-05 

m3120 132 1331 1372 0 nenh l=2e-06 w=4e-06 

m3121 1372 1329 1371 0 nenh l=2e-06 w=4e-06 

m3122 1372 83 1373 0 nenh l=2e-06 w=4e-06 

m3123 1373 81 1374 0 nenh l=2e-06 w=4e-06 

m3124 1374 1375 0 0 nenh l=2e-06 w=4e-06 

m3125 0 1373 1376 0 nenh l=2e-06 w=8e-06 

m3126 1376 74 1375 0 nenh l=2e-06 w=8e-06 

m3127 1371 1375 0 0 nenh l=2e-06 w=4e-06 

m3128 0 1370 731 0 nenh l=2e-06 w=1.4e-05 

m3129 731 1370 0 0 nenh l=2e-06 w=1.9e-05 

m3130 132 1329 1372 3 penh l=2e-06 w=6e-06 

m3131 1372 1331 1371 3 penh l=2e-06 w=6e-06 

m3132 1372 81 1373 3 penh l=2e-06 w=6e-06 

m3133 1373 83 1377 3 penh l=2e-06 w=6e-06 

m3134 1377 1375 3 3 penh l=2e-06 w=6e-06 

m3135 3 1373 1375 3 penh l=2e-06 w=6e-06 

m3136 1375 74 3 3 penh l=2e-06 w=6e-06 

m3137 3 1375 1371 3 penh l=2e-06 w=6e-06 

m3138 3 1371 1370 3 penh l=2e-06 w=2.4e-05 

m3139 3 1370 731 3 penh l=2e-06 w=1.8e-05 

m3140 731 1370 3 3 penh l=2e-06 w=3e-05 

m3141 3 1370 731 3 penh l=2e-06 w=1.8e-05 

m3142 731 1370 3 3 penh l=2e-06 w=2.8e-05 

m3143 139 1329 1378 3 penh l=2e-06 w=6e-06 

m3144 1378 1331 1379 3 penh l=2e-06 w=6e-06 

m3145 1378 81 1380 3 penh l=2e-06 w=6e-06 

m3146 1380 83 1381 3 penh l=2e-06 w=6e-06 

m3147 1381 1382 3 3 penh l=2e-06 w=6e-06 

m3148 3 1380 1382 3 penh l=2e-06 w=6e-06 

m3149 1382 74 3 3 penh l=2e-06 w=6e-06 

m3150 3 1382 1379 3 penh l=2e-06 w=6e-06 

m3151 3 1379 1383 3 penh l=2e-06 w=2.4e-05 

m3152 139 1331 1378 0 nenh l=2e-06 w=4e-06 

m3153 1378 1329 1379 0 nenh l=2e-06 w=4e-06 

m3154 3 1383 697 3 penh l=2e-06 w=2.8e-05 

m3155 697 1383 3 3 penh l=2e-06 w=3e-05 

m3156 697 1383 3 3 penh l=2e-06 w=1.8e-05 

m3157 1378 83 1380 0 nenh l=2e-06 w=4e-06 

m3158 1380 81 1384 0 nenh l=2e-06 w=4e-06 

m3159 1384 1382 0 0 nenh l=2e-06 w=4e-06 

m3160 0 1380 1385 0 nenh l=2e-06 w=8e-06 

m3161 1385 74 1382 0 nenh l=2e-06 w=8e-06 

m3162 3 1383 697 3 penh l=2e-06 w=1.8e-05 

m3163 1379 1382 0 0 nenh l=2e-06 w=4e-06 

m3164 0 1379 1383 0 nenh l=2e-06 w=1.6e-05 

m3165 697 1383 0 0 nenh l=2e-06 w=1.4e-05 

m3166 0 1383 697 0 nenh l=2e-06 w=3.1e-05 

m3167 697 1383 0 0 nenh l=2e-06 w=1.9e-05 

m3168 0 1387 1386 0 nenh l=2e-06 w=1.6e-05 

m3169 0 1386 694 0 nenh l=2e-06 w=3.1e-05 

m3170 152 1331 1388 0 nenh l=2e-06 w=4e-06 

m3171 1388 1329 1387 0 nenh l=2e-06 w=4e-06 

m3172 1388 83 1389 0 nenh l=2e-06 w=4e-06 

m3173 1389 81 1390 0 nenh l=2e-06 w=4e-06 

m3174 1390 1391 0 0 nenh l=2e-06 w=4e-06 

m3175 0 1389 1392 0 nenh l=2e-06 w=8e-06 

m3176 1392 74 1391 0 nenh l=2e-06 w=8e-06 

m3177 1387 1391 0 0 nenh l=2e-06 w=4e-06 

m3178 0 1386 694 0 nenh l=2e-06 w=1.4e-05 

m3179 694 1386 0 0 nenh l=2e-06 w=1.9e-05 

m3180 152 1329 1388 3 penh l=2e-06 w=6e-06 

m3181 1388 1331 1387 3 penh l=2e-06 w=6e-06 

m3182 1388 81 1389 3 penh l=2e-06 w=6e-06 

m3183 1389 83 1393 3 penh l=2e-06 w=6e-06 

m3184 1393 1391 3 3 penh l=2e-06 w=6e-06 

m3185 3 1389 1391 3 penh l=2e-06 w=6e-06 

m3186 1391 74 3 3 penh l=2e-06 w=6e-06 

m3187 3 1391 1387 3 penh l=2e-06 w=6e-06 

m3188 3 1387 1386 3 penh l=2e-06 w=2.4e-05 

m3189 3 1386 694 3 penh l=2e-06 w=1.8e-05 

m3190 694 1386 3 3 penh l=2e-06 w=3e-05 

m3191 3 1386 694 3 penh l=2e-06 w=1.8e-05 

m3192 694 1386 3 3 penh l=2e-06 w=2.8e-05 

m3193 159 1329 1394 3 penh l=2e-06 w=6e-06 

m3194 1394 1331 1395 3 penh l=2e-06 w=6e-06 

m3195 1394 81 1396 3 penh l=2e-06 w=6e-06 

m3196 1396 83 1397 3 penh l=2e-06 w=6e-06 

m3197 1397 1398 3 3 penh l=2e-06 w=6e-06 

m3198 3 1396 1398 3 penh l=2e-06 w=6e-06 

m3199 1398 74 3 3 penh l=2e-06 w=6e-06 

m3200 3 1398 1395 3 penh l=2e-06 w=6e-06 

m3201 3 1395 1399 3 penh l=2e-06 w=2.4e-05 

m3202 159 1331 1394 0 nenh l=2e-06 w=4e-06 

m3203 1394 1329 1395 0 nenh l=2e-06 w=4e-06 

m3204 3 1399 660 3 penh l=2e-06 w=2.8e-05 

m3205 660 1399 3 3 penh l=2e-06 w=3e-05 

m3206 660 1399 3 3 penh l=2e-06 w=1.8e-05 

m3207 1394 83 1396 0 nenh l=2e-06 w=4e-06 

m3208 1396 81 1400 0 nenh l=2e-06 w=4e-06 

m3209 1400 1398 0 0 nenh l=2e-06 w=4e-06 

m3210 0 1396 1401 0 nenh l=2e-06 w=8e-06 

m3211 1401 74 1398 0 nenh l=2e-06 w=8e-06 

m3212 3 1399 660 3 penh l=2e-06 w=1.8e-05 

m3213 1395 1398 0 0 nenh l=2e-06 w=4e-06 

m3214 0 1395 1399 0 nenh l=2e-06 w=1.6e-05 

m3215 660 1399 0 0 nenh l=2e-06 w=1.4e-05 

m3216 0 1399 660 0 nenh l=2e-06 w=3.1e-05 

m3217 660 1399 0 0 nenh l=2e-06 w=1.9e-05 

m3218 0 1403 1402 0 nenh l=2e-06 w=1.6e-05 

m3219 0 1402 657 0 nenh l=2e-06 w=3.1e-05 

m3220 53 1331 1404 0 nenh l=2e-06 w=4e-06 

m3221 1404 1329 1403 0 nenh l=2e-06 w=4e-06 

m3222 1404 83 1405 0 nenh l=2e-06 w=4e-06 

m3223 1405 81 1406 0 nenh l=2e-06 w=4e-06 

m3224 1406 1407 0 0 nenh l=2e-06 w=4e-06 

m3225 0 1405 1408 0 nenh l=2e-06 w=8e-06 

m3226 1408 74 1407 0 nenh l=2e-06 w=8e-06 

m3227 1403 1407 0 0 nenh l=2e-06 w=4e-06 

m3228 0 1402 657 0 nenh l=2e-06 w=1.4e-05 

m3229 657 1402 0 0 nenh l=2e-06 w=1.9e-05 

m3230 53 1329 1404 3 penh l=2e-06 w=6e-06 

m3231 1404 1331 1403 3 penh l=2e-06 w=6e-06 

m3232 1404 81 1405 3 penh l=2e-06 w=6e-06 

m3233 1405 83 1409 3 penh l=2e-06 w=6e-06 

m3234 1409 1407 3 3 penh l=2e-06 w=6e-06 

m3235 3 1405 1407 3 penh l=2e-06 w=6e-06 

m3236 1407 74 3 3 penh l=2e-06 w=6e-06 

m3237 3 1407 1403 3 penh l=2e-06 w=6e-06 

m3238 3 1403 1402 3 penh l=2e-06 w=2.4e-05 

m3239 3 1402 657 3 penh l=2e-06 w=1.8e-05 

m3240 657 1402 3 3 penh l=2e-06 w=3e-05 

m3241 3 1402 657 3 penh l=2e-06 w=1.8e-05 

m3242 657 1402 3 3 penh l=2e-06 w=2.8e-05 

m3243 178 1329 1410 3 penh l=2e-06 w=6e-06 

m3244 1410 1331 1411 3 penh l=2e-06 w=6e-06 

m3245 1410 81 1412 3 penh l=2e-06 w=6e-06 

m3246 1412 83 1413 3 penh l=2e-06 w=6e-06 

m3247 1413 1414 3 3 penh l=2e-06 w=6e-06 

m3248 3 1412 1414 3 penh l=2e-06 w=6e-06 

m3249 1414 74 3 3 penh l=2e-06 w=6e-06 

m3250 3 1414 1411 3 penh l=2e-06 w=6e-06 

m3251 3 1411 1415 3 penh l=2e-06 w=2.4e-05 

m3252 178 1331 1410 0 nenh l=2e-06 w=4e-06 

m3253 1410 1329 1411 0 nenh l=2e-06 w=4e-06 

m3254 3 1415 623 3 penh l=2e-06 w=2.8e-05 

m3255 623 1415 3 3 penh l=2e-06 w=3e-05 

m3256 623 1415 3 3 penh l=2e-06 w=1.8e-05 

m3257 1410 83 1412 0 nenh l=2e-06 w=4e-06 

m3258 1412 81 1416 0 nenh l=2e-06 w=4e-06 

m3259 1416 1414 0 0 nenh l=2e-06 w=4e-06 

m3260 0 1412 1417 0 nenh l=2e-06 w=8e-06 

m3261 1417 74 1414 0 nenh l=2e-06 w=8e-06 

m3262 3 1415 623 3 penh l=2e-06 w=1.8e-05 

m3263 1411 1414 0 0 nenh l=2e-06 w=4e-06 

m3264 0 1411 1415 0 nenh l=2e-06 w=1.6e-05 

m3265 623 1415 0 0 nenh l=2e-06 w=1.4e-05 

m3266 0 1415 623 0 nenh l=2e-06 w=3.1e-05 

m3267 623 1415 0 0 nenh l=2e-06 w=1.9e-05 

m3268 0 1419 1418 0 nenh l=2e-06 w=1.6e-05 

m3269 0 1418 620 0 nenh l=2e-06 w=3.1e-05 

m3270 48 1331 1420 0 nenh l=2e-06 w=4e-06 

m3271 1420 1329 1419 0 nenh l=2e-06 w=4e-06 

m3272 1420 83 1421 0 nenh l=2e-06 w=4e-06 

m3273 1421 81 1422 0 nenh l=2e-06 w=4e-06 

m3274 1422 1423 0 0 nenh l=2e-06 w=4e-06 

m3275 0 1421 1424 0 nenh l=2e-06 w=8e-06 

m3276 1424 74 1423 0 nenh l=2e-06 w=8e-06 

m3277 1419 1423 0 0 nenh l=2e-06 w=4e-06 

m3278 0 1418 620 0 nenh l=2e-06 w=1.4e-05 

m3279 620 1418 0 0 nenh l=2e-06 w=1.9e-05 

m3280 48 1329 1420 3 penh l=2e-06 w=6e-06 

m3281 1420 1331 1419 3 penh l=2e-06 w=6e-06 

m3282 1420 81 1421 3 penh l=2e-06 w=6e-06 

m3283 1421 83 1425 3 penh l=2e-06 w=6e-06 

m3284 1425 1423 3 3 penh l=2e-06 w=6e-06 

m3285 3 1421 1423 3 penh l=2e-06 w=6e-06 

m3286 1423 74 3 3 penh l=2e-06 w=6e-06 

m3287 3 1423 1419 3 penh l=2e-06 w=6e-06 

m3288 3 1419 1418 3 penh l=2e-06 w=2.4e-05 

m3289 3 1418 620 3 penh l=2e-06 w=1.8e-05 

m3290 620 1418 3 3 penh l=2e-06 w=3e-05 

m3291 3 1418 620 3 penh l=2e-06 w=1.8e-05 

m3292 620 1418 3 3 penh l=2e-06 w=2.8e-05 

m3293 197 1329 1426 3 penh l=2e-06 w=6e-06 

m3294 1426 1331 1427 3 penh l=2e-06 w=6e-06 

m3295 1426 81 1428 3 penh l=2e-06 w=6e-06 

m3296 1428 83 1429 3 penh l=2e-06 w=6e-06 

m3297 1429 1430 3 3 penh l=2e-06 w=6e-06 

m3298 3 1428 1430 3 penh l=2e-06 w=6e-06 

m3299 1430 74 3 3 penh l=2e-06 w=6e-06 

m3300 3 1430 1427 3 penh l=2e-06 w=6e-06 

m3301 3 1427 1431 3 penh l=2e-06 w=2.4e-05 

m3302 197 1331 1426 0 nenh l=2e-06 w=4e-06 

m3303 1426 1329 1427 0 nenh l=2e-06 w=4e-06 

m3304 3 1431 586 3 penh l=2e-06 w=2.8e-05 

m3305 586 1431 3 3 penh l=2e-06 w=3e-05 

m3306 586 1431 3 3 penh l=2e-06 w=1.8e-05 

m3307 1426 83 1428 0 nenh l=2e-06 w=4e-06 

m3308 1428 81 1432 0 nenh l=2e-06 w=4e-06 

m3309 1432 1430 0 0 nenh l=2e-06 w=4e-06 

m3310 0 1428 1433 0 nenh l=2e-06 w=8e-06 

m3311 1433 74 1430 0 nenh l=2e-06 w=8e-06 

m3312 3 1431 586 3 penh l=2e-06 w=1.8e-05 

m3313 1427 1430 0 0 nenh l=2e-06 w=4e-06 

m3314 0 1427 1431 0 nenh l=2e-06 w=1.6e-05 

m3315 586 1431 0 0 nenh l=2e-06 w=1.4e-05 

m3316 0 1431 586 0 nenh l=2e-06 w=3.1e-05 

m3317 586 1431 0 0 nenh l=2e-06 w=1.9e-05 

m3318 0 1435 1434 0 nenh l=2e-06 w=1.6e-05 

m3319 0 1434 583 0 nenh l=2e-06 w=3.1e-05 

m3320 43 1331 1436 0 nenh l=2e-06 w=4e-06 

m3321 1436 1329 1435 0 nenh l=2e-06 w=4e-06 

m3322 1436 83 1437 0 nenh l=2e-06 w=4e-06 

m3323 1437 81 1438 0 nenh l=2e-06 w=4e-06 

m3324 1438 1439 0 0 nenh l=2e-06 w=4e-06 

m3325 0 1437 1440 0 nenh l=2e-06 w=8e-06 

m3326 1440 74 1439 0 nenh l=2e-06 w=8e-06 

m3327 1435 1439 0 0 nenh l=2e-06 w=4e-06 

m3328 0 1434 583 0 nenh l=2e-06 w=1.4e-05 

m3329 583 1434 0 0 nenh l=2e-06 w=1.9e-05 

m3330 43 1329 1436 3 penh l=2e-06 w=6e-06 

m3331 1436 1331 1435 3 penh l=2e-06 w=6e-06 

m3332 1436 81 1437 3 penh l=2e-06 w=6e-06 

m3333 1437 83 1441 3 penh l=2e-06 w=6e-06 

m3334 1441 1439 3 3 penh l=2e-06 w=6e-06 

m3335 3 1437 1439 3 penh l=2e-06 w=6e-06 

m3336 1439 74 3 3 penh l=2e-06 w=6e-06 

m3337 3 1439 1435 3 penh l=2e-06 w=6e-06 

m3338 3 1435 1434 3 penh l=2e-06 w=2.4e-05 

m3339 3 1434 583 3 penh l=2e-06 w=1.8e-05 

m3340 583 1434 3 3 penh l=2e-06 w=3e-05 

m3341 3 1434 583 3 penh l=2e-06 w=1.8e-05 

m3342 583 1434 3 3 penh l=2e-06 w=2.8e-05 

m3343 216 1329 1442 3 penh l=2e-06 w=6e-06 

m3344 1442 1331 1443 3 penh l=2e-06 w=6e-06 

m3345 1442 81 1444 3 penh l=2e-06 w=6e-06 

m3346 1444 83 1445 3 penh l=2e-06 w=6e-06 

m3347 1445 1446 3 3 penh l=2e-06 w=6e-06 

m3348 3 1444 1446 3 penh l=2e-06 w=6e-06 

m3349 1446 74 3 3 penh l=2e-06 w=6e-06 

m3350 3 1446 1443 3 penh l=2e-06 w=6e-06 

m3351 3 1443 1447 3 penh l=2e-06 w=2.4e-05 

m3352 216 1331 1442 0 nenh l=2e-06 w=4e-06 

m3353 1442 1329 1443 0 nenh l=2e-06 w=4e-06 

m3354 3 1447 549 3 penh l=2e-06 w=2.8e-05 

m3355 549 1447 3 3 penh l=2e-06 w=3e-05 

m3356 549 1447 3 3 penh l=2e-06 w=1.8e-05 

m3357 1442 83 1444 0 nenh l=2e-06 w=4e-06 

m3358 1444 81 1448 0 nenh l=2e-06 w=4e-06 

m3359 1448 1446 0 0 nenh l=2e-06 w=4e-06 

m3360 0 1444 1449 0 nenh l=2e-06 w=8e-06 

m3361 1449 74 1446 0 nenh l=2e-06 w=8e-06 

m3362 3 1447 549 3 penh l=2e-06 w=1.8e-05 

m3363 1443 1446 0 0 nenh l=2e-06 w=4e-06 

m3364 0 1443 1447 0 nenh l=2e-06 w=1.6e-05 

m3365 549 1447 0 0 nenh l=2e-06 w=1.4e-05 

m3366 0 1447 549 0 nenh l=2e-06 w=3.1e-05 

m3367 549 1447 0 0 nenh l=2e-06 w=1.9e-05 

m3368 0 1451 1450 0 nenh l=2e-06 w=1.6e-05 

m3369 0 1450 546 0 nenh l=2e-06 w=3.1e-05 

m3370 38 1331 1452 0 nenh l=2e-06 w=4e-06 

m3371 1452 1329 1451 0 nenh l=2e-06 w=4e-06 

m3372 1452 83 1453 0 nenh l=2e-06 w=4e-06 

m3373 1453 81 1454 0 nenh l=2e-06 w=4e-06 

m3374 1454 1455 0 0 nenh l=2e-06 w=4e-06 

m3375 0 1453 1456 0 nenh l=2e-06 w=8e-06 

m3376 1456 74 1455 0 nenh l=2e-06 w=8e-06 

m3377 1451 1455 0 0 nenh l=2e-06 w=4e-06 

m3378 0 1450 546 0 nenh l=2e-06 w=1.4e-05 

m3379 546 1450 0 0 nenh l=2e-06 w=1.9e-05 

m3380 38 1329 1452 3 penh l=2e-06 w=6e-06 

m3381 1452 1331 1451 3 penh l=2e-06 w=6e-06 

m3382 1452 81 1453 3 penh l=2e-06 w=6e-06 

m3383 1453 83 1457 3 penh l=2e-06 w=6e-06 

m3384 1457 1455 3 3 penh l=2e-06 w=6e-06 

m3385 3 1453 1455 3 penh l=2e-06 w=6e-06 

m3386 1455 74 3 3 penh l=2e-06 w=6e-06 

m3387 3 1455 1451 3 penh l=2e-06 w=6e-06 

m3388 3 1451 1450 3 penh l=2e-06 w=2.4e-05 

m3389 3 1450 546 3 penh l=2e-06 w=1.8e-05 

m3390 546 1450 3 3 penh l=2e-06 w=3e-05 

m3391 3 1450 546 3 penh l=2e-06 w=1.8e-05 

m3392 546 1450 3 3 penh l=2e-06 w=2.8e-05 

m3393 92 1458 3 3 penh l=2e-06 w=6.2e-05 

m3394 3 1459 1458 3 penh l=2e-06 w=6.2e-05 

m3395 1459 1460 3 3 penh l=2e-06 w=2.9e-05 

m3396 3 1461 1460 3 penh l=4e-06 w=2.9e-05 

m3397 1459 1460 0 0 nenh l=2e-06 w=2.1e-05 

m3398 0 1461 1460 0 nenh l=4e-06 w=2.1e-05 

m3399 92 1458 0 0 nenh l=2e-06 w=4.8e-05 

m3400 0 1459 1458 0 nenh l=2e-06 w=4.8e-05 

m3401 1461 0 0 0 nenh l=4e-06 w=2.5e-05 

m3402 3 1462 79 3 penh l=2e-06 w=5.7e-05 

m3403 3 1463 77 3 penh l=2e-06 w=5.7e-05 

m3404 3 1465 1464 3 penh l=2e-06 w=3.3e-05 

m3405 1464 1466 1463 3 penh l=2e-06 w=3e-05 

m3406 3 1465 1467 3 penh l=2e-06 w=1.5e-05 

m3407 3 1466 1467 3 penh l=2e-06 w=1.5e-05 

m3408 0 1462 79 0 nenh l=2e-06 w=3e-05 

m3409 0 1463 77 0 nenh l=2e-06 w=3e-05 

m3410 3 1467 1331 3 penh l=2e-06 w=5.7e-05 

m3411 3 1468 1462 3 penh l=2e-06 w=1.5e-05 

m3412 3 1469 1462 3 penh l=2e-06 w=1.5e-05 

m3413 0 1465 1463 0 nenh l=2e-06 w=7e-06 

m3414 1463 1466 0 0 nenh l=2e-06 w=7e-06 

m3415 3 1468 1466 3 penh l=2e-06 w=1.3e-05 

m3416 3 1469 1470 3 penh l=2e-06 w=3.3e-05 

m3417 1470 1466 1471 3 penh l=2e-06 w=3e-05 

m3418 1472 1465 0 0 nenh l=2e-06 w=1.6e-05 

m3419 1472 1466 1467 0 nenh l=2e-06 w=1.4e-05 

m3420 0 1467 1331 0 nenh l=2e-06 w=3e-05 

m3421 3 1473 1329 3 penh l=2e-06 w=5.7e-05 

m3422 3 1468 1474 3 penh l=2e-06 w=3.3e-05 

m3423 1474 1469 1473 3 penh l=2e-06 w=3e-05 

m3424 3 1465 1475 3 penh l=2e-06 w=1.5e-05 

m3425 3 1465 1469 3 penh l=2e-06 w=1.3e-05 

m3426 3 1468 1475 3 penh l=2e-06 w=1.5e-05 

m3427 1476 1468 0 0 nenh l=2e-06 w=1.6e-05 

m3428 1476 1469 1462 0 nenh l=2e-06 w=1.4e-05 

m3429 0 1468 1466 0 nenh l=2e-06 w=7e-06 

m3430 0 1469 1471 0 nenh l=2e-06 w=7e-06 

m3431 1471 1466 0 0 nenh l=2e-06 w=7e-06 

m3432 0 1473 1329 0 nenh l=2e-06 w=3e-05 

m3433 3 1471 1477 3 penh l=2e-06 w=5.7e-05 

m3434 0 1468 1473 0 nenh l=2e-06 w=7e-06 

m3435 1473 1469 0 0 nenh l=2e-06 w=7e-06 

m3436 0 1465 1469 0 nenh l=2e-06 w=7e-06 

m3437 3 1475 1478 3 penh l=2e-06 w=5.7e-05 

m3438 1479 1465 0 0 nenh l=2e-06 w=1.6e-05 

m3439 1479 1468 1475 0 nenh l=2e-06 w=1.4e-05 

m3440 0 1471 1477 0 nenh l=2e-06 w=3e-05 

m3441 0 1475 1478 0 nenh l=2e-06 w=3e-05 

m3442 1468 1480 3 3 penh l=2e-06 w=6.2e-05 

m3443 3 1481 1480 3 penh l=2e-06 w=6.2e-05 

m3444 1481 1482 3 3 penh l=2e-06 w=2.9e-05 

m3445 3 1483 1482 3 penh l=4e-06 w=2.9e-05 

m3446 1481 1482 0 0 nenh l=2e-06 w=2.1e-05 

m3447 0 1483 1482 0 nenh l=4e-06 w=2.1e-05 

m3448 1468 1480 0 0 nenh l=2e-06 w=4.8e-05 

m3449 0 1481 1480 0 nenh l=2e-06 w=4.8e-05 

m3450 1483 0 0 0 nenh l=4e-06 w=2.5e-05 

m3451 1465 1484 3 3 penh l=2e-06 w=6.2e-05 

m3452 3 1485 1484 3 penh l=2e-06 w=6.2e-05 

m3453 1485 1486 3 3 penh l=2e-06 w=2.9e-05 

m3454 3 1487 1486 3 penh l=4e-06 w=2.9e-05 

m3455 1485 1486 0 0 nenh l=2e-06 w=2.1e-05 

m3456 0 1487 1486 0 nenh l=4e-06 w=2.1e-05 

m3457 1465 1484 0 0 nenh l=2e-06 w=4.8e-05 

m3458 0 1485 1484 0 nenh l=2e-06 w=4.8e-05 

m3459 1487 0 0 0 nenh l=4e-06 w=2.5e-05 

m3460 75 1488 3 3 penh l=2e-06 w=6.2e-05 

m3461 3 1489 1488 3 penh l=2e-06 w=6.2e-05 

m3462 1489 1490 3 3 penh l=2e-06 w=2.9e-05 

m3463 3 1491 1490 3 penh l=4e-06 w=2.9e-05 

m3464 1489 1490 0 0 nenh l=2e-06 w=2.1e-05 

m3465 0 1491 1490 0 nenh l=4e-06 w=2.1e-05 

m3466 75 1488 0 0 nenh l=2e-06 w=4.8e-05 

m3467 0 1489 1488 0 nenh l=2e-06 w=4.8e-05 

m3468 1491 0 0 0 nenh l=4e-06 w=2.5e-05 

m3469 99 1492 3 3 penh l=2e-06 w=6.2e-05 

m3470 3 1493 1492 3 penh l=2e-06 w=6.2e-05 

m3471 1493 1494 3 3 penh l=2e-06 w=2.9e-05 

m3472 3 1495 1494 3 penh l=4e-06 w=2.9e-05 

m3473 1493 1494 0 0 nenh l=2e-06 w=2.1e-05 

m3474 0 1495 1494 0 nenh l=4e-06 w=2.1e-05 

m3475 99 1492 0 0 nenh l=2e-06 w=4.8e-05 

m3476 0 1493 1492 0 nenh l=2e-06 w=4.8e-05 

m3477 1495 0 0 0 nenh l=4e-06 w=2.5e-05 

m3478 3 1497 1496 3 penh l=2e-06 w=9.7e-05 

m3479 1496 1497 3 3 penh l=2e-06 w=9.5e-05 

m3480 3 1497 1496 3 penh l=2e-06 w=9.5e-05 

m3481 1496 1497 3 3 penh l=2e-06 w=9.6e-05 

m3482 3 1497 1496 3 penh l=2e-06 w=9.6e-05 

m3483 1496 1497 3 3 penh l=2e-06 w=9.5e-05 

m3484 3 1497 1496 3 penh l=2e-06 w=9.5e-05 

m3485 1496 1497 3 3 penh l=2e-06 w=9.6e-05 

m3486 3 1498 1497 3 penh l=2e-06 w=5.3e-05 

m3487 1497 1498 3 3 penh l=2e-06 w=5.3e-05 

m3488 3 1499 1498 3 penh l=2e-06 w=4.9e-05 

m3489 1499 282 3 3 penh l=2e-06 w=2.3e-05 

m3490 3 1498 1497 3 penh l=2e-06 w=4.8e-05 

m3491 1497 1498 3 3 penh l=2e-06 w=4.8e-05 

m3492 3 282 1500 3 penh l=2e-06 w=2.2e-05 

m3493 1501 1502 3 3 penh l=2e-06 w=5e-05 

m3494 3 1500 1502 3 penh l=2e-06 w=4.7e-05 

m3495 1501 1502 3 3 penh l=2e-06 w=4.8e-05 

m3496 3 1502 1501 3 penh l=2e-06 w=4.8e-05 

m3497 0 1501 1496 0 nenh l=2e-06 w=4.6e-05 

m3498 1496 1501 0 0 nenh l=2e-06 w=4.8e-05 

m3499 0 1501 1496 0 nenh l=2e-06 w=4.6e-05 

m3500 1496 1501 0 0 nenh l=2e-06 w=4.8e-05 

m3501 0 1501 1496 0 nenh l=2e-06 w=4.8e-05 

m3502 1496 1501 0 0 nenh l=2e-06 w=4.8e-05 

m3503 0 1501 1496 0 nenh l=2e-06 w=4.8e-05 

m3504 1496 1501 0 0 nenh l=2e-06 w=4.6e-05 

m3505 0 1502 1501 0 nenh l=2e-06 w=6e-05 

m3506 1501 1502 0 0 nenh l=2e-06 w=6e-05 

m3507 1502 1500 0 0 nenh l=2e-06 w=5e-05 

m3508 0 1498 1497 0 nenh l=2e-06 w=3.5e-05 

m3509 1497 1498 0 0 nenh l=2e-06 w=3.4e-05 

m3510 0 282 1500 0 nenh l=2e-06 w=2.4e-05 

m3511 0 1498 1497 0 nenh l=2e-06 w=2.5e-05 

m3512 1497 1498 0 0 nenh l=2e-06 w=2.5e-05 

m3513 0 1499 1498 0 nenh l=2e-06 w=1.6e-05 

m3514 1499 282 0 0 nenh l=2e-06 w=2.3e-05 

m3515 3 1503 327 3 penh l=2e-06 w=0.0001 

m3516 327 1503 3 3 penh l=2e-06 w=0.0001 

m3517 3 1503 327 3 penh l=2e-06 w=0.0001 

m3518 327 1503 3 3 penh l=2e-06 w=0.0001 

m3519 3 1503 327 3 penh l=2e-06 w=0.0001 

m3520 327 1503 3 3 penh l=2e-06 w=0.0001 

m3521 3 1503 327 3 penh l=2e-06 w=0.0001 

m3522 327 1503 3 3 penh l=2e-06 w=0.0001 

m3523 0 1503 327 0 nenh l=2e-06 w=9.7e-05 

m3524 327 1503 0 0 nenh l=2e-06 w=9.7e-05 

m3525 0 1503 327 0 nenh l=2e-06 w=9.7e-05 

m3526 327 1503 0 0 nenh l=2e-06 w=9.7e-05 

m3527 3 1504 329 3 penh l=2e-06 w=0.0001 

m3528 329 1504 3 3 penh l=2e-06 w=0.0001 

m3529 3 1504 329 3 penh l=2e-06 w=0.0001 

m3530 329 1504 3 3 penh l=2e-06 w=0.0001 

m3531 3 1504 329 3 penh l=2e-06 w=0.0001 

m3532 329 1504 3 3 penh l=2e-06 w=0.0001 

m3533 3 1504 329 3 penh l=2e-06 w=0.0001 

m3534 329 1504 3 3 penh l=2e-06 w=0.0001 

m3535 0 1504 329 0 nenh l=2e-06 w=9.7e-05 

m3536 329 1504 0 0 nenh l=2e-06 w=9.7e-05 

m3537 0 1504 329 0 nenh l=2e-06 w=9.7e-05 

m3538 329 1504 0 0 nenh l=2e-06 w=9.7e-05 

m3539 3 1505 81 3 penh l=2e-06 w=0.0001 

m3540 81 1505 3 3 penh l=2e-06 w=0.0001 

m3541 3 1505 81 3 penh l=2e-06 w=0.0001 

m3542 81 1505 3 3 penh l=2e-06 w=0.0001 

m3543 3 1505 81 3 penh l=2e-06 w=0.0001 

m3544 81 1505 3 3 penh l=2e-06 w=0.0001 

m3545 3 1505 81 3 penh l=2e-06 w=0.0001 

m3546 81 1505 3 3 penh l=2e-06 w=0.0001 

m3547 0 1505 81 0 nenh l=2e-06 w=9.7e-05 

m3548 81 1505 0 0 nenh l=2e-06 w=9.7e-05 

m3549 0 1505 81 0 nenh l=2e-06 w=9.7e-05 

m3550 81 1505 0 0 nenh l=2e-06 w=9.7e-05 

m3551 3 1506 83 3 penh l=2e-06 w=0.0001 

m3552 83 1506 3 3 penh l=2e-06 w=0.0001 

m3553 3 1506 83 3 penh l=2e-06 w=0.0001 

m3554 83 1506 3 3 penh l=2e-06 w=0.0001 

m3555 3 1506 83 3 penh l=2e-06 w=0.0001 

m3556 83 1506 3 3 penh l=2e-06 w=0.0001 

m3557 3 1506 83 3 penh l=2e-06 w=0.0001 

m3558 83 1506 3 3 penh l=2e-06 w=0.0001 

m3559 0 1506 83 0 nenh l=2e-06 w=9.7e-05 

m3560 83 1506 0 0 nenh l=2e-06 w=9.7e-05 

m3561 0 1506 83 0 nenh l=2e-06 w=9.7e-05 

m3562 83 1506 0 0 nenh l=2e-06 w=9.7e-05 

m3563 0 1507 1506 0 nenh l=2e-06 w=2.9e-05 

m3564 1506 1507 0 0 nenh l=2e-06 w=1.7e-05 

m3565 0 1507 1506 0 nenh l=2e-06 w=2.9e-05 

m3566 1506 1507 0 0 nenh l=2e-06 w=1.7e-05 

m3567 0 1507 1506 0 nenh l=2e-06 w=1.2e-05 

m3568 0 1508 1504 0 nenh l=2e-06 w=2.9e-05 

m3569 1504 1508 0 0 nenh l=2e-06 w=1.7e-05 

m3570 0 1507 1506 0 nenh l=2e-06 w=1.2e-05 

m3571 0 1508 1504 0 nenh l=2e-06 w=2.9e-05 

m3572 1504 1508 0 0 nenh l=2e-06 w=1.7e-05 

m3573 0 1508 1504 0 nenh l=2e-06 w=1.2e-05 

m3574 0 1508 1504 0 nenh l=2e-06 w=1.2e-05 

m3575 1506 1507 3 3 penh l=2e-06 w=2.2e-05 

m3576 3 1507 1506 3 penh l=2e-06 w=3.4e-05 

m3577 1506 1507 3 3 penh l=2e-06 w=2.3e-05 

m3578 1506 1507 3 3 penh l=2e-06 w=2.2e-05 

m3579 3 1507 1506 3 penh l=2e-06 w=3.4e-05 

m3580 1506 1507 3 3 penh l=2e-06 w=2.3e-05 

m3581 1509 81 0 0 nenh l=2e-06 w=1.4e-05 

m3582 0 1510 1503 0 nenh l=2e-06 w=2.9e-05 

m3583 0 83 1511 0 nenh l=2e-06 w=7e-06 

m3584 1511 1509 0 0 nenh l=2e-06 w=7e-06 

m3585 0 1512 1511 0 nenh l=2e-06 w=7e-06 

m3586 1504 1508 3 3 penh l=2e-06 w=2.2e-05 

m3587 3 1508 1504 3 penh l=2e-06 w=3.4e-05 

m3588 1504 1508 3 3 penh l=2e-06 w=2.3e-05 

m3589 1504 1508 3 3 penh l=2e-06 w=2.2e-05 

m3590 3 1508 1504 3 penh l=2e-06 w=3.4e-05 

m3591 1504 1508 3 3 penh l=2e-06 w=2.3e-05 

m3592 0 1511 1510 0 nenh l=2e-06 w=3e-05 

m3593 1503 1510 0 0 nenh l=2e-06 w=1.7e-05 

m3594 0 1510 1503 0 nenh l=2e-06 w=2.9e-05 

m3595 1503 1510 0 0 nenh l=2e-06 w=1.7e-05 

m3596 0 1510 1503 0 nenh l=2e-06 w=1.2e-05 

m3597 0 1510 1503 0 nenh l=2e-06 w=1.2e-05 

m3598 1513 83 1511 3 penh l=2e-06 w=3.4e-05 

m3599 1506 1507 3 3 penh l=2e-06 w=2.7e-05 

m3600 1506 1507 3 3 penh l=2e-06 w=2.7e-05 

m3601 1504 1508 3 3 penh l=2e-06 w=2.7e-05 

m3602 1504 1508 3 3 penh l=2e-06 w=2.7e-05 

m3603 1509 81 3 3 penh l=2e-06 w=3.1e-05 

m3604 1513 1509 1514 3 penh l=2e-06 w=3.4e-05 

m3605 1514 1512 3 3 penh l=2e-06 w=3.5e-05 

m3606 3 1511 1510 3 penh l=2e-06 w=5.7e-05 

m3607 1515 329 0 0 nenh l=2e-06 w=1.4e-05 

m3608 1503 1510 3 3 penh l=2e-06 w=2.2e-05 

m3609 3 1510 1503 3 penh l=2e-06 w=3.4e-05 

m3610 1503 1510 3 3 penh l=2e-06 w=2.3e-05 

m3611 1503 1510 3 3 penh l=2e-06 w=2.2e-05 

m3612 3 1510 1503 3 penh l=2e-06 w=3.4e-05 

m3613 1503 1510 3 3 penh l=2e-06 w=2.3e-05 

m3614 1503 1510 3 3 penh l=2e-06 w=2.7e-05 

m3615 1503 1510 3 3 penh l=2e-06 w=2.7e-05 

m3616 1515 329 3 3 penh l=2e-06 w=3.1e-05 

m3617 0 1516 1505 0 nenh l=2e-06 w=2.9e-05 

m3618 1505 1516 0 0 nenh l=2e-06 w=1.7e-05 

m3619 0 1516 1505 0 nenh l=2e-06 w=2.9e-05 

m3620 1505 1516 0 0 nenh l=2e-06 w=1.7e-05 

m3621 0 1516 1505 0 nenh l=2e-06 w=1.2e-05 

m3622 0 1516 1505 0 nenh l=2e-06 w=1.2e-05 

m3623 0 1517 1508 0 nenh l=2e-06 w=3e-05 

m3624 1518 81 1517 0 nenh l=2e-06 w=1.9e-05 

m3625 1505 1516 3 3 penh l=2e-06 w=2.2e-05 

m3626 3 1516 1505 3 penh l=2e-06 w=3.4e-05 

m3627 1505 1516 3 3 penh l=2e-06 w=2.3e-05 

m3628 1505 1516 3 3 penh l=2e-06 w=2.2e-05 

m3629 3 1516 1505 3 penh l=2e-06 w=3.4e-05 

m3630 1505 1516 3 3 penh l=2e-06 w=2.3e-05 

m3631 1518 1520 1519 0 nenh l=2e-06 w=2e-05 

m3632 1519 1521 0 0 nenh l=2e-06 w=2.6e-05 

m3633 1520 83 0 0 nenh l=2e-06 w=1.4e-05 

m3634 0 1522 1516 0 nenh l=2e-06 w=3e-05 

m3635 1521 1512 0 0 nenh l=2e-06 w=1.4e-05 

m3636 0 329 1522 0 nenh l=2e-06 w=7e-06 

m3637 1522 1523 0 0 nenh l=2e-06 w=7e-06 

m3638 0 1521 1522 0 nenh l=2e-06 w=7e-06 

m3639 1505 1516 3 3 penh l=2e-06 w=2.7e-05 

m3640 1505 1516 3 3 penh l=2e-06 w=2.7e-05 

m3641 3 1517 1508 3 penh l=2e-06 w=5.7e-05 

m3642 1520 83 3 3 penh l=2e-06 w=3.1e-05 

m3643 1517 81 3 3 penh l=2e-06 w=1.4e-05 

m3644 3 1520 1517 3 penh l=2e-06 w=1.5e-05 

m3645 1517 1521 3 3 penh l=2e-06 w=1.7e-05 

m3646 3 1522 1516 3 penh l=2e-06 w=5.7e-05 

m3647 0 1524 1507 0 nenh l=2e-06 w=3e-05 

m3648 1523 327 0 0 nenh l=2e-06 w=1.4e-05 

m3649 1525 327 1524 0 nenh l=2e-06 w=1.9e-05 

m3650 1526 329 1522 3 penh l=2e-06 w=3.4e-05 

m3651 1521 1512 3 3 penh l=2e-06 w=3.1e-05 

m3652 1526 1523 1527 3 penh l=2e-06 w=3.4e-05 

m3653 1527 1521 3 3 penh l=2e-06 w=3.5e-05 

m3654 3 1524 1507 3 penh l=2e-06 w=5.7e-05 

m3655 1525 1515 1528 0 nenh l=2e-06 w=2e-05 

m3656 1528 1512 0 0 nenh l=2e-06 w=2.6e-05 

m3657 1523 327 3 3 penh l=2e-06 w=3.1e-05 

m3658 1524 327 3 3 penh l=2e-06 w=1.4e-05 

m3659 3 1515 1524 3 penh l=2e-06 w=1.5e-05 

m3660 1524 1512 3 3 penh l=2e-06 w=1.7e-05 

m3661 75 1477 1529 3 penh l=2e-06 w=6e-06 

m3662 1529 1478 1530 3 penh l=2e-06 w=6e-06 

m3663 1529 81 1531 3 penh l=2e-06 w=6e-06 

m3664 1531 83 1532 3 penh l=2e-06 w=6e-06 

m3665 1532 1533 3 3 penh l=2e-06 w=6e-06 

m3666 3 1531 1533 3 penh l=2e-06 w=6e-06 

m3667 1533 74 3 3 penh l=2e-06 w=6e-06 

m3668 3 1533 1530 3 penh l=2e-06 w=6e-06 

m3669 3 1530 1534 3 penh l=2e-06 w=2.4e-05 

m3670 75 1478 1529 0 nenh l=2e-06 w=4e-06 

m3671 1529 1477 1530 0 nenh l=2e-06 w=4e-06 

m3672 3 1534 810 3 penh l=2e-06 w=2.8e-05 

m3673 810 1534 3 3 penh l=2e-06 w=3e-05 

m3674 810 1534 3 3 penh l=2e-06 w=1.8e-05 

m3675 1529 83 1531 0 nenh l=2e-06 w=4e-06 

m3676 1531 81 1535 0 nenh l=2e-06 w=4e-06 

m3677 1535 1533 0 0 nenh l=2e-06 w=4e-06 

m3678 0 1531 1536 0 nenh l=2e-06 w=8e-06 

m3679 1536 74 1533 0 nenh l=2e-06 w=8e-06 

m3680 3 1534 810 3 penh l=2e-06 w=1.8e-05 

m3681 1530 1533 0 0 nenh l=2e-06 w=4e-06 

m3682 0 1530 1534 0 nenh l=2e-06 w=1.6e-05 

m3683 810 1534 0 0 nenh l=2e-06 w=1.4e-05 

m3684 0 1534 810 0 nenh l=2e-06 w=3.1e-05 

m3685 810 1534 0 0 nenh l=2e-06 w=1.9e-05 

m3686 0 1538 1537 0 nenh l=2e-06 w=1.6e-05 

m3687 0 1537 803 0 nenh l=2e-06 w=3.1e-05 

m3688 92 1478 1539 0 nenh l=2e-06 w=4e-06 

m3689 1539 1477 1538 0 nenh l=2e-06 w=4e-06 

m3690 1539 83 1540 0 nenh l=2e-06 w=4e-06 

m3691 1540 81 1541 0 nenh l=2e-06 w=4e-06 

m3692 1541 1542 0 0 nenh l=2e-06 w=4e-06 

m3693 0 1540 1543 0 nenh l=2e-06 w=8e-06 

m3694 1543 74 1542 0 nenh l=2e-06 w=8e-06 

m3695 1538 1542 0 0 nenh l=2e-06 w=4e-06 

m3696 0 1537 803 0 nenh l=2e-06 w=1.4e-05 

m3697 803 1537 0 0 nenh l=2e-06 w=1.9e-05 

m3698 92 1477 1539 3 penh l=2e-06 w=6e-06 

m3699 1539 1478 1538 3 penh l=2e-06 w=6e-06 

m3700 1539 81 1540 3 penh l=2e-06 w=6e-06 

m3701 1540 83 1544 3 penh l=2e-06 w=6e-06 

m3702 1544 1542 3 3 penh l=2e-06 w=6e-06 

m3703 3 1540 1542 3 penh l=2e-06 w=6e-06 

m3704 1542 74 3 3 penh l=2e-06 w=6e-06 

m3705 3 1542 1538 3 penh l=2e-06 w=6e-06 

m3706 3 1538 1537 3 penh l=2e-06 w=2.4e-05 

m3707 3 1537 803 3 penh l=2e-06 w=1.8e-05 

m3708 803 1537 3 3 penh l=2e-06 w=3e-05 

m3709 3 1537 803 3 penh l=2e-06 w=1.8e-05 

m3710 803 1537 3 3 penh l=2e-06 w=2.8e-05 

m3711 99 1477 1545 3 penh l=2e-06 w=6e-06 

m3712 1545 1478 1546 3 penh l=2e-06 w=6e-06 

m3713 1545 81 1547 3 penh l=2e-06 w=6e-06 

m3714 1547 83 1548 3 penh l=2e-06 w=6e-06 

m3715 1548 1549 3 3 penh l=2e-06 w=6e-06 

m3716 3 1547 1549 3 penh l=2e-06 w=6e-06 

m3717 1549 74 3 3 penh l=2e-06 w=6e-06 

m3718 3 1549 1546 3 penh l=2e-06 w=6e-06 

m3719 3 1546 1550 3 penh l=2e-06 w=2.4e-05 

m3720 99 1478 1545 0 nenh l=2e-06 w=4e-06 

m3721 1545 1477 1546 0 nenh l=2e-06 w=4e-06 

m3722 3 1550 773 3 penh l=2e-06 w=2.8e-05 

m3723 773 1550 3 3 penh l=2e-06 w=3e-05 

m3724 773 1550 3 3 penh l=2e-06 w=1.8e-05 

m3725 1545 83 1547 0 nenh l=2e-06 w=4e-06 

m3726 1547 81 1551 0 nenh l=2e-06 w=4e-06 

m3727 1551 1549 0 0 nenh l=2e-06 w=4e-06 

m3728 0 1547 1552 0 nenh l=2e-06 w=8e-06 

m3729 1552 74 1549 0 nenh l=2e-06 w=8e-06 

m3730 3 1550 773 3 penh l=2e-06 w=1.8e-05 

m3731 1546 1549 0 0 nenh l=2e-06 w=4e-06 

m3732 0 1546 1550 0 nenh l=2e-06 w=1.6e-05 

m3733 773 1550 0 0 nenh l=2e-06 w=1.4e-05 

m3734 0 1550 773 0 nenh l=2e-06 w=3.1e-05 

m3735 773 1550 0 0 nenh l=2e-06 w=1.9e-05 

m3736 0 1554 1553 0 nenh l=2e-06 w=1.6e-05 

m3737 0 1553 766 0 nenh l=2e-06 w=3.1e-05 

m3738 112 1478 1555 0 nenh l=2e-06 w=4e-06 

m3739 1555 1477 1554 0 nenh l=2e-06 w=4e-06 

m3740 1555 83 1556 0 nenh l=2e-06 w=4e-06 

m3741 1556 81 1557 0 nenh l=2e-06 w=4e-06 

m3742 1557 1558 0 0 nenh l=2e-06 w=4e-06 

m3743 0 1556 1559 0 nenh l=2e-06 w=8e-06 

m3744 1559 74 1558 0 nenh l=2e-06 w=8e-06 

m3745 1554 1558 0 0 nenh l=2e-06 w=4e-06 

m3746 0 1553 766 0 nenh l=2e-06 w=1.4e-05 

m3747 766 1553 0 0 nenh l=2e-06 w=1.9e-05 

m3748 112 1477 1555 3 penh l=2e-06 w=6e-06 

m3749 1555 1478 1554 3 penh l=2e-06 w=6e-06 

m3750 1555 81 1556 3 penh l=2e-06 w=6e-06 

m3751 1556 83 1560 3 penh l=2e-06 w=6e-06 

m3752 1560 1558 3 3 penh l=2e-06 w=6e-06 

m3753 3 1556 1558 3 penh l=2e-06 w=6e-06 

m3754 1558 74 3 3 penh l=2e-06 w=6e-06 

m3755 3 1558 1554 3 penh l=2e-06 w=6e-06 

m3756 3 1554 1553 3 penh l=2e-06 w=2.4e-05 

m3757 3 1553 766 3 penh l=2e-06 w=1.8e-05 

m3758 766 1553 3 3 penh l=2e-06 w=3e-05 

m3759 3 1553 766 3 penh l=2e-06 w=1.8e-05 

m3760 766 1553 3 3 penh l=2e-06 w=2.8e-05 

m3761 119 1477 1561 3 penh l=2e-06 w=6e-06 

m3762 1561 1478 1562 3 penh l=2e-06 w=6e-06 

m3763 1561 81 1563 3 penh l=2e-06 w=6e-06 

m3764 1563 83 1564 3 penh l=2e-06 w=6e-06 

m3765 1564 1565 3 3 penh l=2e-06 w=6e-06 

m3766 3 1563 1565 3 penh l=2e-06 w=6e-06 

m3767 1565 74 3 3 penh l=2e-06 w=6e-06 

m3768 3 1565 1562 3 penh l=2e-06 w=6e-06 

m3769 3 1562 1566 3 penh l=2e-06 w=2.4e-05 

m3770 119 1478 1561 0 nenh l=2e-06 w=4e-06 

m3771 1561 1477 1562 0 nenh l=2e-06 w=4e-06 

m3772 3 1566 736 3 penh l=2e-06 w=2.8e-05 

m3773 736 1566 3 3 penh l=2e-06 w=3e-05 

m3774 736 1566 3 3 penh l=2e-06 w=1.8e-05 

m3775 1561 83 1563 0 nenh l=2e-06 w=4e-06 

m3776 1563 81 1567 0 nenh l=2e-06 w=4e-06 

m3777 1567 1565 0 0 nenh l=2e-06 w=4e-06 

m3778 0 1563 1568 0 nenh l=2e-06 w=8e-06 

m3779 1568 74 1565 0 nenh l=2e-06 w=8e-06 

m3780 3 1566 736 3 penh l=2e-06 w=1.8e-05 

m3781 1562 1565 0 0 nenh l=2e-06 w=4e-06 

m3782 0 1562 1566 0 nenh l=2e-06 w=1.6e-05 

m3783 736 1566 0 0 nenh l=2e-06 w=1.4e-05 

m3784 0 1566 736 0 nenh l=2e-06 w=3.1e-05 

m3785 736 1566 0 0 nenh l=2e-06 w=1.9e-05 

m3786 0 1570 1569 0 nenh l=2e-06 w=1.6e-05 

m3787 0 1569 729 0 nenh l=2e-06 w=3.1e-05 

m3788 132 1478 1571 0 nenh l=2e-06 w=4e-06 

m3789 1571 1477 1570 0 nenh l=2e-06 w=4e-06 

m3790 1571 83 1572 0 nenh l=2e-06 w=4e-06 

m3791 1572 81 1573 0 nenh l=2e-06 w=4e-06 

m3792 1573 1574 0 0 nenh l=2e-06 w=4e-06 

m3793 0 1572 1575 0 nenh l=2e-06 w=8e-06 

m3794 1575 74 1574 0 nenh l=2e-06 w=8e-06 

m3795 1570 1574 0 0 nenh l=2e-06 w=4e-06 

m3796 0 1569 729 0 nenh l=2e-06 w=1.4e-05 

m3797 729 1569 0 0 nenh l=2e-06 w=1.9e-05 

m3798 132 1477 1571 3 penh l=2e-06 w=6e-06 

m3799 1571 1478 1570 3 penh l=2e-06 w=6e-06 

m3800 1571 81 1572 3 penh l=2e-06 w=6e-06 

m3801 1572 83 1576 3 penh l=2e-06 w=6e-06 

m3802 1576 1574 3 3 penh l=2e-06 w=6e-06 

m3803 3 1572 1574 3 penh l=2e-06 w=6e-06 

m3804 1574 74 3 3 penh l=2e-06 w=6e-06 

m3805 3 1574 1570 3 penh l=2e-06 w=6e-06 

m3806 3 1570 1569 3 penh l=2e-06 w=2.4e-05 

m3807 3 1569 729 3 penh l=2e-06 w=1.8e-05 

m3808 729 1569 3 3 penh l=2e-06 w=3e-05 

m3809 3 1569 729 3 penh l=2e-06 w=1.8e-05 

m3810 729 1569 3 3 penh l=2e-06 w=2.8e-05 

m3811 139 1477 1577 3 penh l=2e-06 w=6e-06 

m3812 1577 1478 1578 3 penh l=2e-06 w=6e-06 

m3813 1577 81 1579 3 penh l=2e-06 w=6e-06 

m3814 1579 83 1580 3 penh l=2e-06 w=6e-06 

m3815 1580 1581 3 3 penh l=2e-06 w=6e-06 

m3816 3 1579 1581 3 penh l=2e-06 w=6e-06 

m3817 1581 74 3 3 penh l=2e-06 w=6e-06 

m3818 3 1581 1578 3 penh l=2e-06 w=6e-06 

m3819 3 1578 1582 3 penh l=2e-06 w=2.4e-05 

m3820 139 1478 1577 0 nenh l=2e-06 w=4e-06 

m3821 1577 1477 1578 0 nenh l=2e-06 w=4e-06 

m3822 3 1582 699 3 penh l=2e-06 w=2.8e-05 

m3823 699 1582 3 3 penh l=2e-06 w=3e-05 

m3824 699 1582 3 3 penh l=2e-06 w=1.8e-05 

m3825 1577 83 1579 0 nenh l=2e-06 w=4e-06 

m3826 1579 81 1583 0 nenh l=2e-06 w=4e-06 

m3827 1583 1581 0 0 nenh l=2e-06 w=4e-06 

m3828 0 1579 1584 0 nenh l=2e-06 w=8e-06 

m3829 1584 74 1581 0 nenh l=2e-06 w=8e-06 

m3830 3 1582 699 3 penh l=2e-06 w=1.8e-05 

m3831 1578 1581 0 0 nenh l=2e-06 w=4e-06 

m3832 0 1578 1582 0 nenh l=2e-06 w=1.6e-05 

m3833 699 1582 0 0 nenh l=2e-06 w=1.4e-05 

m3834 0 1582 699 0 nenh l=2e-06 w=3.1e-05 

m3835 699 1582 0 0 nenh l=2e-06 w=1.9e-05 

m3836 0 1586 1585 0 nenh l=2e-06 w=1.6e-05 

m3837 0 1585 692 0 nenh l=2e-06 w=3.1e-05 

m3838 152 1478 1587 0 nenh l=2e-06 w=4e-06 

m3839 1587 1477 1586 0 nenh l=2e-06 w=4e-06 

m3840 1587 83 1588 0 nenh l=2e-06 w=4e-06 

m3841 1588 81 1589 0 nenh l=2e-06 w=4e-06 

m3842 1589 1590 0 0 nenh l=2e-06 w=4e-06 

m3843 0 1588 1591 0 nenh l=2e-06 w=8e-06 

m3844 1591 74 1590 0 nenh l=2e-06 w=8e-06 

m3845 1586 1590 0 0 nenh l=2e-06 w=4e-06 

m3846 0 1585 692 0 nenh l=2e-06 w=1.4e-05 

m3847 692 1585 0 0 nenh l=2e-06 w=1.9e-05 

m3848 152 1477 1587 3 penh l=2e-06 w=6e-06 

m3849 1587 1478 1586 3 penh l=2e-06 w=6e-06 

m3850 1587 81 1588 3 penh l=2e-06 w=6e-06 

m3851 1588 83 1592 3 penh l=2e-06 w=6e-06 

m3852 1592 1590 3 3 penh l=2e-06 w=6e-06 

m3853 3 1588 1590 3 penh l=2e-06 w=6e-06 

m3854 1590 74 3 3 penh l=2e-06 w=6e-06 

m3855 3 1590 1586 3 penh l=2e-06 w=6e-06 

m3856 3 1586 1585 3 penh l=2e-06 w=2.4e-05 

m3857 3 1585 692 3 penh l=2e-06 w=1.8e-05 

m3858 692 1585 3 3 penh l=2e-06 w=3e-05 

m3859 3 1585 692 3 penh l=2e-06 w=1.8e-05 

m3860 692 1585 3 3 penh l=2e-06 w=2.8e-05 

m3861 159 1477 1593 3 penh l=2e-06 w=6e-06 

m3862 1593 1478 1594 3 penh l=2e-06 w=6e-06 

m3863 1593 81 1595 3 penh l=2e-06 w=6e-06 

m3864 1595 83 1596 3 penh l=2e-06 w=6e-06 

m3865 1596 1597 3 3 penh l=2e-06 w=6e-06 

m3866 3 1595 1597 3 penh l=2e-06 w=6e-06 

m3867 1597 74 3 3 penh l=2e-06 w=6e-06 

m3868 3 1597 1594 3 penh l=2e-06 w=6e-06 

m3869 3 1594 1598 3 penh l=2e-06 w=2.4e-05 

m3870 159 1478 1593 0 nenh l=2e-06 w=4e-06 

m3871 1593 1477 1594 0 nenh l=2e-06 w=4e-06 

m3872 3 1598 662 3 penh l=2e-06 w=2.8e-05 

m3873 662 1598 3 3 penh l=2e-06 w=3e-05 

m3874 662 1598 3 3 penh l=2e-06 w=1.8e-05 

m3875 1593 83 1595 0 nenh l=2e-06 w=4e-06 

m3876 1595 81 1599 0 nenh l=2e-06 w=4e-06 

m3877 1599 1597 0 0 nenh l=2e-06 w=4e-06 

m3878 0 1595 1600 0 nenh l=2e-06 w=8e-06 

m3879 1600 74 1597 0 nenh l=2e-06 w=8e-06 

m3880 3 1598 662 3 penh l=2e-06 w=1.8e-05 

m3881 1594 1597 0 0 nenh l=2e-06 w=4e-06 

m3882 0 1594 1598 0 nenh l=2e-06 w=1.6e-05 

m3883 662 1598 0 0 nenh l=2e-06 w=1.4e-05 

m3884 0 1598 662 0 nenh l=2e-06 w=3.1e-05 

m3885 662 1598 0 0 nenh l=2e-06 w=1.9e-05 

m3886 0 1602 1601 0 nenh l=2e-06 w=1.6e-05 

m3887 0 1601 655 0 nenh l=2e-06 w=3.1e-05 

m3888 53 1478 1603 0 nenh l=2e-06 w=4e-06 

m3889 1603 1477 1602 0 nenh l=2e-06 w=4e-06 

m3890 1603 83 1604 0 nenh l=2e-06 w=4e-06 

m3891 1604 81 1605 0 nenh l=2e-06 w=4e-06 

m3892 1605 1606 0 0 nenh l=2e-06 w=4e-06 

m3893 0 1604 1607 0 nenh l=2e-06 w=8e-06 

m3894 1607 74 1606 0 nenh l=2e-06 w=8e-06 

m3895 1602 1606 0 0 nenh l=2e-06 w=4e-06 

m3896 0 1601 655 0 nenh l=2e-06 w=1.4e-05 

m3897 655 1601 0 0 nenh l=2e-06 w=1.9e-05 

m3898 53 1477 1603 3 penh l=2e-06 w=6e-06 

m3899 1603 1478 1602 3 penh l=2e-06 w=6e-06 

m3900 1603 81 1604 3 penh l=2e-06 w=6e-06 

m3901 1604 83 1608 3 penh l=2e-06 w=6e-06 

m3902 1608 1606 3 3 penh l=2e-06 w=6e-06 

m3903 3 1604 1606 3 penh l=2e-06 w=6e-06 

m3904 1606 74 3 3 penh l=2e-06 w=6e-06 

m3905 3 1606 1602 3 penh l=2e-06 w=6e-06 

m3906 3 1602 1601 3 penh l=2e-06 w=2.4e-05 

m3907 3 1601 655 3 penh l=2e-06 w=1.8e-05 

m3908 655 1601 3 3 penh l=2e-06 w=3e-05 

m3909 3 1601 655 3 penh l=2e-06 w=1.8e-05 

m3910 655 1601 3 3 penh l=2e-06 w=2.8e-05 

m3911 178 1477 1609 3 penh l=2e-06 w=6e-06 

m3912 1609 1478 1610 3 penh l=2e-06 w=6e-06 

m3913 1609 81 1611 3 penh l=2e-06 w=6e-06 

m3914 1611 83 1612 3 penh l=2e-06 w=6e-06 

m3915 1612 1613 3 3 penh l=2e-06 w=6e-06 

m3916 3 1611 1613 3 penh l=2e-06 w=6e-06 

m3917 1613 74 3 3 penh l=2e-06 w=6e-06 

m3918 3 1613 1610 3 penh l=2e-06 w=6e-06 

m3919 3 1610 1614 3 penh l=2e-06 w=2.4e-05 

m3920 178 1478 1609 0 nenh l=2e-06 w=4e-06 

m3921 1609 1477 1610 0 nenh l=2e-06 w=4e-06 

m3922 3 1614 625 3 penh l=2e-06 w=2.8e-05 

m3923 625 1614 3 3 penh l=2e-06 w=3e-05 

m3924 625 1614 3 3 penh l=2e-06 w=1.8e-05 

m3925 1609 83 1611 0 nenh l=2e-06 w=4e-06 

m3926 1611 81 1615 0 nenh l=2e-06 w=4e-06 

m3927 1615 1613 0 0 nenh l=2e-06 w=4e-06 

m3928 0 1611 1616 0 nenh l=2e-06 w=8e-06 

m3929 1616 74 1613 0 nenh l=2e-06 w=8e-06 

m3930 3 1614 625 3 penh l=2e-06 w=1.8e-05 

m3931 1610 1613 0 0 nenh l=2e-06 w=4e-06 

m3932 0 1610 1614 0 nenh l=2e-06 w=1.6e-05 

m3933 625 1614 0 0 nenh l=2e-06 w=1.4e-05 

m3934 0 1614 625 0 nenh l=2e-06 w=3.1e-05 

m3935 625 1614 0 0 nenh l=2e-06 w=1.9e-05 

m3936 0 1618 1617 0 nenh l=2e-06 w=1.6e-05 

m3937 0 1617 618 0 nenh l=2e-06 w=3.1e-05 

m3938 48 1478 1619 0 nenh l=2e-06 w=4e-06 

m3939 1619 1477 1618 0 nenh l=2e-06 w=4e-06 

m3940 1619 83 1620 0 nenh l=2e-06 w=4e-06 

m3941 1620 81 1621 0 nenh l=2e-06 w=4e-06 

m3942 1621 1622 0 0 nenh l=2e-06 w=4e-06 

m3943 0 1620 1623 0 nenh l=2e-06 w=8e-06 

m3944 1623 74 1622 0 nenh l=2e-06 w=8e-06 

m3945 1618 1622 0 0 nenh l=2e-06 w=4e-06 

m3946 0 1617 618 0 nenh l=2e-06 w=1.4e-05 

m3947 618 1617 0 0 nenh l=2e-06 w=1.9e-05 

m3948 48 1477 1619 3 penh l=2e-06 w=6e-06 

m3949 1619 1478 1618 3 penh l=2e-06 w=6e-06 

m3950 1619 81 1620 3 penh l=2e-06 w=6e-06 

m3951 1620 83 1624 3 penh l=2e-06 w=6e-06 

m3952 1624 1622 3 3 penh l=2e-06 w=6e-06 

m3953 3 1620 1622 3 penh l=2e-06 w=6e-06 

m3954 1622 74 3 3 penh l=2e-06 w=6e-06 

m3955 3 1622 1618 3 penh l=2e-06 w=6e-06 

m3956 3 1618 1617 3 penh l=2e-06 w=2.4e-05 

m3957 3 1617 618 3 penh l=2e-06 w=1.8e-05 

m3958 618 1617 3 3 penh l=2e-06 w=3e-05 

m3959 3 1617 618 3 penh l=2e-06 w=1.8e-05 

m3960 618 1617 3 3 penh l=2e-06 w=2.8e-05 

m3961 197 1477 1625 3 penh l=2e-06 w=6e-06 

m3962 1625 1478 1626 3 penh l=2e-06 w=6e-06 

m3963 1625 81 1627 3 penh l=2e-06 w=6e-06 

m3964 1627 83 1628 3 penh l=2e-06 w=6e-06 

m3965 1628 1629 3 3 penh l=2e-06 w=6e-06 

m3966 3 1627 1629 3 penh l=2e-06 w=6e-06 

m3967 1629 74 3 3 penh l=2e-06 w=6e-06 

m3968 3 1629 1626 3 penh l=2e-06 w=6e-06 

m3969 3 1626 1630 3 penh l=2e-06 w=2.4e-05 

m3970 197 1478 1625 0 nenh l=2e-06 w=4e-06 

m3971 1625 1477 1626 0 nenh l=2e-06 w=4e-06 

m3972 3 1630 588 3 penh l=2e-06 w=2.8e-05 

m3973 588 1630 3 3 penh l=2e-06 w=3e-05 

m3974 588 1630 3 3 penh l=2e-06 w=1.8e-05 

m3975 1625 83 1627 0 nenh l=2e-06 w=4e-06 

m3976 1627 81 1631 0 nenh l=2e-06 w=4e-06 

m3977 1631 1629 0 0 nenh l=2e-06 w=4e-06 

m3978 0 1627 1632 0 nenh l=2e-06 w=8e-06 

m3979 1632 74 1629 0 nenh l=2e-06 w=8e-06 

m3980 3 1630 588 3 penh l=2e-06 w=1.8e-05 

m3981 1626 1629 0 0 nenh l=2e-06 w=4e-06 

m3982 0 1626 1630 0 nenh l=2e-06 w=1.6e-05 

m3983 588 1630 0 0 nenh l=2e-06 w=1.4e-05 

m3984 0 1630 588 0 nenh l=2e-06 w=3.1e-05 

m3985 588 1630 0 0 nenh l=2e-06 w=1.9e-05 

m3986 0 1634 1633 0 nenh l=2e-06 w=1.6e-05 

m3987 0 1633 581 0 nenh l=2e-06 w=3.1e-05 

m3988 43 1478 1635 0 nenh l=2e-06 w=4e-06 

m3989 1635 1477 1634 0 nenh l=2e-06 w=4e-06 

m3990 1635 83 1636 0 nenh l=2e-06 w=4e-06 

m3991 1636 81 1637 0 nenh l=2e-06 w=4e-06 

m3992 1637 1638 0 0 nenh l=2e-06 w=4e-06 

m3993 0 1636 1639 0 nenh l=2e-06 w=8e-06 

m3994 1639 74 1638 0 nenh l=2e-06 w=8e-06 

m3995 1634 1638 0 0 nenh l=2e-06 w=4e-06 

m3996 0 1633 581 0 nenh l=2e-06 w=1.4e-05 

m3997 581 1633 0 0 nenh l=2e-06 w=1.9e-05 

m3998 43 1477 1635 3 penh l=2e-06 w=6e-06 

m3999 1635 1478 1634 3 penh l=2e-06 w=6e-06 

m4000 1635 81 1636 3 penh l=2e-06 w=6e-06 

m4001 1636 83 1640 3 penh l=2e-06 w=6e-06 

m4002 1640 1638 3 3 penh l=2e-06 w=6e-06 

m4003 3 1636 1638 3 penh l=2e-06 w=6e-06 

m4004 1638 74 3 3 penh l=2e-06 w=6e-06 

m4005 3 1638 1634 3 penh l=2e-06 w=6e-06 

m4006 3 1634 1633 3 penh l=2e-06 w=2.4e-05 

m4007 3 1633 581 3 penh l=2e-06 w=1.8e-05 

m4008 581 1633 3 3 penh l=2e-06 w=3e-05 

m4009 3 1633 581 3 penh l=2e-06 w=1.8e-05 

m4010 581 1633 3 3 penh l=2e-06 w=2.8e-05 

m4011 216 1477 1641 3 penh l=2e-06 w=6e-06 

m4012 1641 1478 1642 3 penh l=2e-06 w=6e-06 

m4013 1641 81 1643 3 penh l=2e-06 w=6e-06 

m4014 1643 83 1644 3 penh l=2e-06 w=6e-06 

m4015 1644 1645 3 3 penh l=2e-06 w=6e-06 

m4016 3 1643 1645 3 penh l=2e-06 w=6e-06 

m4017 1645 74 3 3 penh l=2e-06 w=6e-06 

m4018 3 1645 1642 3 penh l=2e-06 w=6e-06 

m4019 3 1642 1646 3 penh l=2e-06 w=2.4e-05 

m4020 216 1478 1641 0 nenh l=2e-06 w=4e-06 

m4021 1641 1477 1642 0 nenh l=2e-06 w=4e-06 

m4022 3 1646 551 3 penh l=2e-06 w=2.8e-05 

m4023 551 1646 3 3 penh l=2e-06 w=3e-05 

m4024 551 1646 3 3 penh l=2e-06 w=1.8e-05 

m4025 1641 83 1643 0 nenh l=2e-06 w=4e-06 

m4026 1643 81 1647 0 nenh l=2e-06 w=4e-06 

m4027 1647 1645 0 0 nenh l=2e-06 w=4e-06 

m4028 0 1643 1648 0 nenh l=2e-06 w=8e-06 

m4029 1648 74 1645 0 nenh l=2e-06 w=8e-06 

m4030 3 1646 551 3 penh l=2e-06 w=1.8e-05 

m4031 1642 1645 0 0 nenh l=2e-06 w=4e-06 

m4032 0 1642 1646 0 nenh l=2e-06 w=1.6e-05 

m4033 551 1646 0 0 nenh l=2e-06 w=1.4e-05 

m4034 0 1646 551 0 nenh l=2e-06 w=3.1e-05 

m4035 551 1646 0 0 nenh l=2e-06 w=1.9e-05 

m4036 0 1650 1649 0 nenh l=2e-06 w=1.6e-05 

m4037 0 1649 544 0 nenh l=2e-06 w=3.1e-05 

m4038 38 1478 1651 0 nenh l=2e-06 w=4e-06 

m4039 1651 1477 1650 0 nenh l=2e-06 w=4e-06 

m4040 1651 83 1652 0 nenh l=2e-06 w=4e-06 

m4041 1652 81 1653 0 nenh l=2e-06 w=4e-06 

m4042 1653 1654 0 0 nenh l=2e-06 w=4e-06 

m4043 0 1652 1655 0 nenh l=2e-06 w=8e-06 

m4044 1655 74 1654 0 nenh l=2e-06 w=8e-06 

m4045 1650 1654 0 0 nenh l=2e-06 w=4e-06 

m4046 0 1649 544 0 nenh l=2e-06 w=1.4e-05 

m4047 544 1649 0 0 nenh l=2e-06 w=1.9e-05 

m4048 38 1477 1651 3 penh l=2e-06 w=6e-06 

m4049 1651 1478 1650 3 penh l=2e-06 w=6e-06 

m4050 1651 81 1652 3 penh l=2e-06 w=6e-06 

m4051 1652 83 1656 3 penh l=2e-06 w=6e-06 

m4052 1656 1654 3 3 penh l=2e-06 w=6e-06 

m4053 3 1652 1654 3 penh l=2e-06 w=6e-06 

m4054 1654 74 3 3 penh l=2e-06 w=6e-06 

m4055 3 1654 1650 3 penh l=2e-06 w=6e-06 

m4056 3 1650 1649 3 penh l=2e-06 w=2.4e-05 

m4057 3 1649 544 3 penh l=2e-06 w=1.8e-05 

m4058 544 1649 3 3 penh l=2e-06 w=3e-05 

m4059 3 1649 544 3 penh l=2e-06 w=1.8e-05 

m4060 544 1649 3 3 penh l=2e-06 w=2.8e-05 

m4061 119 1657 3 3 penh l=2e-06 w=6.2e-05 

m4062 3 1658 1657 3 penh l=2e-06 w=6.2e-05 

m4063 1658 1659 3 3 penh l=2e-06 w=2.9e-05 

m4064 3 1660 1659 3 penh l=4e-06 w=2.9e-05 

m4065 1658 1659 0 0 nenh l=2e-06 w=2.1e-05 

m4066 0 1660 1659 0 nenh l=4e-06 w=2.1e-05 

m4067 119 1657 0 0 nenh l=2e-06 w=4.8e-05 

m4068 0 1658 1657 0 nenh l=2e-06 w=4.8e-05 

m4069 1660 0 0 0 nenh l=4e-06 w=2.5e-05 

m4070 139 1661 3 3 penh l=2e-06 w=6.2e-05 

m4071 3 1662 1661 3 penh l=2e-06 w=6.2e-05 

m4072 1662 1663 3 3 penh l=2e-06 w=2.9e-05 

m4073 3 1664 1663 3 penh l=4e-06 w=2.9e-05 

m4074 1662 1663 0 0 nenh l=2e-06 w=2.1e-05 

m4075 0 1664 1663 0 nenh l=4e-06 w=2.1e-05 

m4076 139 1661 0 0 nenh l=2e-06 w=4.8e-05 

m4077 0 1662 1661 0 nenh l=2e-06 w=4.8e-05 

m4078 1664 0 0 0 nenh l=4e-06 w=2.5e-05 

m4079 3 1666 1665 3 penh l=2e-06 w=9.7e-05 

m4080 1665 1666 3 3 penh l=2e-06 w=9.5e-05 

m4081 3 1666 1665 3 penh l=2e-06 w=9.5e-05 

m4082 1665 1666 3 3 penh l=2e-06 w=9.6e-05 

m4083 3 1666 1665 3 penh l=2e-06 w=9.6e-05 

m4084 1665 1666 3 3 penh l=2e-06 w=9.5e-05 

m4085 3 1666 1665 3 penh l=2e-06 w=9.5e-05 

m4086 1665 1666 3 3 penh l=2e-06 w=9.6e-05 

m4087 3 1667 1666 3 penh l=2e-06 w=5.3e-05 

m4088 1666 1667 3 3 penh l=2e-06 w=5.3e-05 

m4089 3 1668 1667 3 penh l=2e-06 w=4.9e-05 

m4090 1668 277 3 3 penh l=2e-06 w=2.3e-05 

m4091 3 1667 1666 3 penh l=2e-06 w=4.8e-05 

m4092 1666 1667 3 3 penh l=2e-06 w=4.8e-05 

m4093 3 277 1669 3 penh l=2e-06 w=2.2e-05 

m4094 1670 1671 3 3 penh l=2e-06 w=5e-05 

m4095 3 1669 1671 3 penh l=2e-06 w=4.7e-05 

m4096 1670 1671 3 3 penh l=2e-06 w=4.8e-05 

m4097 3 1671 1670 3 penh l=2e-06 w=4.8e-05 

m4098 0 1670 1665 0 nenh l=2e-06 w=4.6e-05 

m4099 1665 1670 0 0 nenh l=2e-06 w=4.8e-05 

m4100 0 1670 1665 0 nenh l=2e-06 w=4.6e-05 

m4101 1665 1670 0 0 nenh l=2e-06 w=4.8e-05 

m4102 0 1670 1665 0 nenh l=2e-06 w=4.8e-05 

m4103 1665 1670 0 0 nenh l=2e-06 w=4.8e-05 

m4104 0 1670 1665 0 nenh l=2e-06 w=4.8e-05 

m4105 1665 1670 0 0 nenh l=2e-06 w=4.6e-05 

m4106 0 1671 1670 0 nenh l=2e-06 w=6e-05 

m4107 1670 1671 0 0 nenh l=2e-06 w=6e-05 

m4108 1671 1669 0 0 nenh l=2e-06 w=5e-05 

m4109 0 1667 1666 0 nenh l=2e-06 w=3.5e-05 

m4110 1666 1667 0 0 nenh l=2e-06 w=3.4e-05 

m4111 0 277 1669 0 nenh l=2e-06 w=2.4e-05 

m4112 0 1667 1666 0 nenh l=2e-06 w=2.5e-05 

m4113 1666 1667 0 0 nenh l=2e-06 w=2.5e-05 

m4114 0 1668 1667 0 nenh l=2e-06 w=1.6e-05 

m4115 1668 277 0 0 nenh l=2e-06 w=2.3e-05 

m4116 857 1672 3 3 penh l=2e-06 w=6.2e-05 

m4117 3 1673 1672 3 penh l=2e-06 w=6.2e-05 

m4118 1673 1674 3 3 penh l=2e-06 w=2.9e-05 

m4119 3 1675 1674 3 penh l=4e-06 w=2.9e-05 

m4120 1673 1674 0 0 nenh l=2e-06 w=2.1e-05 

m4121 0 1675 1674 0 nenh l=4e-06 w=2.1e-05 

m4122 857 1672 0 0 nenh l=2e-06 w=4.8e-05 

m4123 0 1673 1672 0 nenh l=2e-06 w=4.8e-05 

m4124 1675 0 0 0 nenh l=4e-06 w=2.5e-05 

m4125 3 1677 1676 3 penh l=2e-06 w=9.7e-05 

m4126 1676 1677 3 3 penh l=2e-06 w=9.5e-05 

m4127 3 1677 1676 3 penh l=2e-06 w=9.5e-05 

m4128 1676 1677 3 3 penh l=2e-06 w=9.6e-05 

m4129 3 1677 1676 3 penh l=2e-06 w=9.6e-05 

m4130 1676 1677 3 3 penh l=2e-06 w=9.5e-05 

m4131 3 1677 1676 3 penh l=2e-06 w=9.5e-05 

m4132 1676 1677 3 3 penh l=2e-06 w=9.6e-05 

m4133 3 1678 1677 3 penh l=2e-06 w=5.3e-05 

m4134 1677 1678 3 3 penh l=2e-06 w=5.3e-05 

m4135 3 1679 1678 3 penh l=2e-06 w=4.9e-05 

m4136 1679 1319 3 3 penh l=2e-06 w=2.3e-05 

m4137 3 1678 1677 3 penh l=2e-06 w=4.8e-05 

m4138 1677 1678 3 3 penh l=2e-06 w=4.8e-05 

m4139 3 1319 1680 3 penh l=2e-06 w=2.2e-05 

m4140 1681 1682 3 3 penh l=2e-06 w=5e-05 

m4141 3 1680 1682 3 penh l=2e-06 w=4.7e-05 

m4142 1681 1682 3 3 penh l=2e-06 w=4.8e-05 

m4143 3 1682 1681 3 penh l=2e-06 w=4.8e-05 

m4144 0 1681 1676 0 nenh l=2e-06 w=4.6e-05 

m4145 1676 1681 0 0 nenh l=2e-06 w=4.8e-05 

m4146 0 1681 1676 0 nenh l=2e-06 w=4.6e-05 

m4147 1676 1681 0 0 nenh l=2e-06 w=4.8e-05 

m4148 0 1681 1676 0 nenh l=2e-06 w=4.8e-05 

m4149 1676 1681 0 0 nenh l=2e-06 w=4.8e-05 

m4150 0 1681 1676 0 nenh l=2e-06 w=4.8e-05 

m4151 1676 1681 0 0 nenh l=2e-06 w=4.6e-05 

m4152 0 1682 1681 0 nenh l=2e-06 w=6e-05 

m4153 1681 1682 0 0 nenh l=2e-06 w=6e-05 

m4154 1682 1680 0 0 nenh l=2e-06 w=5e-05 

m4155 0 1678 1677 0 nenh l=2e-06 w=3.5e-05 

m4156 1677 1678 0 0 nenh l=2e-06 w=3.4e-05 

m4157 0 1319 1680 0 nenh l=2e-06 w=2.4e-05 

m4158 0 1678 1677 0 nenh l=2e-06 w=2.5e-05 

m4159 1677 1678 0 0 nenh l=2e-06 w=2.5e-05 

m4160 0 1679 1678 0 nenh l=2e-06 w=1.6e-05 

m4161 1679 1319 0 0 nenh l=2e-06 w=2.3e-05 

m4162 1512 1683 3 3 penh l=2e-06 w=6.2e-05 

m4163 3 1684 1683 3 penh l=2e-06 w=6.2e-05 

m4164 1684 1685 3 3 penh l=2e-06 w=2.9e-05 

m4165 3 1686 1685 3 penh l=4e-06 w=2.9e-05 

m4166 1684 1685 0 0 nenh l=2e-06 w=2.1e-05 

m4167 0 1686 1685 0 nenh l=4e-06 w=2.1e-05 

m4168 1512 1683 0 0 nenh l=2e-06 w=4.8e-05 

m4169 0 1684 1683 0 nenh l=2e-06 w=4.8e-05 

m4170 1686 0 0 0 nenh l=4e-06 w=2.5e-05 

m4171 3 1688 1687 3 penh l=2e-06 w=9.7e-05 

m4172 1687 1688 3 3 penh l=2e-06 w=9.5e-05 

m4173 3 1688 1687 3 penh l=2e-06 w=9.5e-05 

m4174 1687 1688 3 3 penh l=2e-06 w=9.6e-05 

m4175 3 1688 1687 3 penh l=2e-06 w=9.6e-05 

m4176 1687 1688 3 3 penh l=2e-06 w=9.5e-05 

m4177 3 1688 1687 3 penh l=2e-06 w=9.5e-05 

m4178 1687 1688 3 3 penh l=2e-06 w=9.6e-05 

m4179 3 1689 1688 3 penh l=2e-06 w=5.3e-05 

m4180 1688 1689 3 3 penh l=2e-06 w=5.3e-05 

m4181 3 1690 1689 3 penh l=2e-06 w=4.9e-05 

m4182 1690 1325 3 3 penh l=2e-06 w=2.3e-05 

m4183 3 1689 1688 3 penh l=2e-06 w=4.8e-05 

m4184 1688 1689 3 3 penh l=2e-06 w=4.8e-05 

m4185 3 1325 1691 3 penh l=2e-06 w=2.2e-05 

m4186 1692 1693 3 3 penh l=2e-06 w=5e-05 

m4187 3 1691 1693 3 penh l=2e-06 w=4.7e-05 

m4188 1692 1693 3 3 penh l=2e-06 w=4.8e-05 

m4189 3 1693 1692 3 penh l=2e-06 w=4.8e-05 

m4190 0 1692 1687 0 nenh l=2e-06 w=4.6e-05 

m4191 1687 1692 0 0 nenh l=2e-06 w=4.8e-05 

m4192 0 1692 1687 0 nenh l=2e-06 w=4.6e-05 

m4193 1687 1692 0 0 nenh l=2e-06 w=4.8e-05 

m4194 0 1692 1687 0 nenh l=2e-06 w=4.8e-05 

m4195 1687 1692 0 0 nenh l=2e-06 w=4.8e-05 

m4196 0 1692 1687 0 nenh l=2e-06 w=4.8e-05 

m4197 1687 1692 0 0 nenh l=2e-06 w=4.6e-05 

m4198 0 1693 1692 0 nenh l=2e-06 w=6e-05 

m4199 1692 1693 0 0 nenh l=2e-06 w=6e-05 

m4200 1693 1691 0 0 nenh l=2e-06 w=5e-05 

m4201 0 1689 1688 0 nenh l=2e-06 w=3.5e-05 

m4202 1688 1689 0 0 nenh l=2e-06 w=3.4e-05 

m4203 0 1325 1691 0 nenh l=2e-06 w=2.4e-05 

m4204 0 1689 1688 0 nenh l=2e-06 w=2.5e-05 

m4205 1688 1689 0 0 nenh l=2e-06 w=2.5e-05 

m4206 0 1690 1689 0 nenh l=2e-06 w=1.6e-05 

m4207 1690 1325 0 0 nenh l=2e-06 w=2.3e-05 

m4208 216 1694 3 3 penh l=2e-06 w=6.2e-05 

m4209 3 1695 1694 3 penh l=2e-06 w=6.2e-05 

m4210 1695 1696 3 3 penh l=2e-06 w=2.9e-05 

m4211 3 1697 1696 3 penh l=4e-06 w=2.9e-05 

m4212 1695 1696 0 0 nenh l=2e-06 w=2.1e-05 

m4213 0 1697 1696 0 nenh l=4e-06 w=2.1e-05 

m4214 216 1694 0 0 nenh l=2e-06 w=4.8e-05 

m4215 0 1695 1694 0 nenh l=2e-06 w=4.8e-05 

m4216 1697 0 0 0 nenh l=4e-06 w=2.5e-05 

m4217 197 1698 3 3 penh l=2e-06 w=6.2e-05 

m4218 3 1699 1698 3 penh l=2e-06 w=6.2e-05 

m4219 1699 1700 3 3 penh l=2e-06 w=2.9e-05 

m4220 3 1701 1700 3 penh l=4e-06 w=2.9e-05 

m4221 1699 1700 0 0 nenh l=2e-06 w=2.1e-05 

m4222 0 1701 1700 0 nenh l=4e-06 w=2.1e-05 

m4223 197 1698 0 0 nenh l=2e-06 w=4.8e-05 

m4224 0 1699 1698 0 nenh l=2e-06 w=4.8e-05 

m4225 1701 0 0 0 nenh l=4e-06 w=2.5e-05 

m4226 178 1702 3 3 penh l=2e-06 w=6.2e-05 

m4227 3 1703 1702 3 penh l=2e-06 w=6.2e-05 

m4228 1703 1704 3 3 penh l=2e-06 w=2.9e-05 

m4229 3 1705 1704 3 penh l=4e-06 w=2.9e-05 

m4230 1703 1704 0 0 nenh l=2e-06 w=2.1e-05 

m4231 0 1705 1704 0 nenh l=4e-06 w=2.1e-05 

m4232 178 1702 0 0 nenh l=2e-06 w=4.8e-05 

m4233 0 1703 1702 0 nenh l=2e-06 w=4.8e-05 

m4234 1705 0 0 0 nenh l=4e-06 w=2.5e-05 

m4235 159 1706 3 3 penh l=2e-06 w=6.2e-05 

m4236 3 1707 1706 3 penh l=2e-06 w=6.2e-05 

m4237 1707 1708 3 3 penh l=2e-06 w=2.9e-05 

m4238 3 1709 1708 3 penh l=4e-06 w=2.9e-05 

m4239 1707 1708 0 0 nenh l=2e-06 w=2.1e-05 

m4240 0 1709 1708 0 nenh l=4e-06 w=2.1e-05 

m4241 159 1706 0 0 nenh l=2e-06 w=4.8e-05 

m4242 0 1707 1706 0 nenh l=2e-06 w=4.8e-05 

m4243 1709 0 0 0 nenh l=4e-06 w=2.5e-05 

c1 21 0 1.38e-13
c2 846 0 1.05e-13
c3 329 0 1.44e-13
c4 57 0 4.1e-13
c5 248 0 1.38e-13
c6 1491 0 4.1e-13
c7 0 0 4.1e-13
c8 0 0 4.1e-13
c9 12 0 1.05e-13
c10 0 0 1.238e-12
c11 1495 0 4.1e-13
c12 847 0 1.38e-13
c13 66 0 1.05e-13
c14 81 0 1.04e-13
c15 329 0 1.99e-13
c16 42 0 4.1e-13
c17 37 0 4.1e-13
c18 263 0 1.05e-13
c19 1461 0 4.1e-13
c20 238 0 4.1e-13
c21 239 0 1.05e-13
c22 327 0 1.24e-13
c23 1487 0 4.1e-13
c24 839 0 1.05e-13
c25 834 0 4.1e-13
c26 67 0 1.38e-13
c27 0 0 4.1e-13
c28 1677 0 1.38e-13
c29 1687 0 1.05e-13
c30 1496 0 1.05e-13
c31 13 0 1.38e-13
c32 47 0 4.1e-13
c33 74 0 1.31e-13
c34 327 0 1.13e-13
c35 255 0 1.05e-13
c36 0 0 4.1e-13
c37 0 0 4.1e-13
c38 840 0 1.38e-13
c39 58 0 1.05e-13
c40 4 0 1.05e-13
c41 3 0 1.05e-13
c42 838 0 4.1e-13
c43 0 0 4.1e-13
c44 1688 0 1.38e-13
c45 1676 0 1.05e-13
c46 74 0 1.32e-13
c47 256 0 1.38e-13
c48 1483 0 4.1e-13
c49 52 0 4.1e-13
c50 20 0 1.05e-13
c51 240 0 1.38e-13
c52 264 0 1.38e-13
c53 59 0 1.38e-13
c54 0 0 4.1e-13
c55 5 0 1.38e-13
c56 3 0 1.38e-13
c57 1497 0 1.38e-13
c58 247 0 1.05e-13
c59 0 0 4.1e-13
c60 32 0 4.1e-13
c61 0 0 9.0322e-11
c67 1709 0 4e-11
c68 1708 0 1.1e-13
c69 159 0 7.01e-13
c70 1707 0 1.15e-13
c71 1706 0 2.2e-13
c72 1705 0 4e-11
c73 1704 0 1.1e-13
c74 178 0 6.92e-13
c75 1703 0 1.15e-13
c76 1702 0 2.2e-13
c77 1701 0 4e-11
c78 1700 0 1.1e-13
c79 197 0 6.82e-13
c80 1699 0 1.15e-13
c81 1698 0 2.2e-13
c82 1697 0 4e-11
c83 1696 0 1.1e-13
c84 216 0 6.66e-13
c85 1695 0 1.15e-13
c86 1694 0 2.2e-13
c87 1692 0 4.38e-13
c88 1693 0 2.03e-13
c89 1691 0 1.23e-13
c90 1325 0 1.66e-13
c91 1690 0 1.21e-13
c92 1689 0 1.91e-13
c93 1687 0 4e-11
c94 1688 0 3.85e-13
c95 1686 0 4e-11
c96 1685 0 1.1e-13
c97 1512 0 2.6e-13
c98 1684 0 1.15e-13
c99 1683 0 2.2e-13
c100 1681 0 4.38e-13
c101 1682 0 2.03e-13
c102 1680 0 1.23e-13
c103 1319 0 2.13e-13
c104 1679 0 1.21e-13
c105 1678 0 1.91e-13
c106 1676 0 4e-11
c107 1677 0 3.85e-13
c108 1675 0 4e-11
c109 1674 0 1.1e-13
c110 857 0 6.72e-13
c111 1673 0 1.15e-13
c112 1672 0 2.2e-13
c113 3 0 1.11603e-10
c114 1670 0 4.38e-13
c115 1671 0 2.03e-13
c116 1669 0 1.23e-13
c117 277 0 1.93e-13
c118 1668 0 1.21e-13
c119 1667 0 1.91e-13
c120 1665 0 4e-11
c121 1666 0 3.85e-13
c123 1664 0 4e-11
c124 1663 0 1.1e-13
c125 1662 0 1.15e-13
c126 1661 0 2.2e-13
c127 1660 0 4e-11
c128 1659 0 1.1e-13
c129 1658 0 1.15e-13
c130 1657 0 2.2e-13
c131 544 0 5.47e-13
c132 551 0 5.51e-13
c133 581 0 5.42e-13
c134 588 0 5.44e-13
c135 618 0 5.41e-13
c136 625 0 5.46e-13
c137 655 0 5.43e-13
c138 662 0 5.44e-13
c139 692 0 5.5e-13
c140 699 0 5.61e-13
c141 729 0 5.48e-13
c142 736 0 5.56e-13
c143 766 0 5.46e-13
c144 773 0 5.43e-13
c145 803 0 5.43e-13
c146 38 0 6.6e-13
c147 43 0 6.69e-13
c148 48 0 6.84e-13
c149 53 0 6.99e-13
c150 152 0 7.2e-13
c151 139 0 7.24e-13
c152 132 0 7.29e-13
c153 119 0 7.37e-13
c154 112 0 7.39e-13
c155 99 0 7.45e-13
c156 92 0 7.46e-13
c157 75 0 7.56e-13
c158 810 0 5.45e-13
c159 1478 0 4.47e-13
c160 1477 0 3.11e-13
c161 74 0 1.336e-12
c162 327 0 2.839e-12
c163 1521 0 1.02e-13
c164 1516 0 1.2e-13
c165 329 0 4.564e-12
c166 1510 0 1.12e-13
c167 1508 0 1.18e-13
c168 1507 0 1.27e-13
c169 83 0 2.978e-12
c170 1506 0 2.93e-13
c171 81 0 2.915e-12
c172 1505 0 2.98e-13
c173 1504 0 3.09e-13
c174 1503 0 3.05e-13
c175 1501 0 4.38e-13
c176 1502 0 2.03e-13
c177 1500 0 1.23e-13
c178 282 0 1.62e-13
c179 1499 0 1.21e-13
c180 1498 0 1.91e-13
c181 1496 0 4e-11
c182 1497 0 3.85e-13
c183 1495 0 4e-11
c184 1494 0 1.1e-13
c185 1493 0 1.15e-13
c186 1492 0 2.2e-13
c187 1491 0 4e-11
c188 1490 0 1.1e-13
c189 1489 0 1.15e-13
c190 1488 0 2.2e-13
c191 1487 0 2.022e-12
c192 1486 0 1.1e-13
c193 1485 0 1.15e-13
c194 1484 0 2.2e-13
c195 1483 0 2.022e-12
c196 1482 0 1.1e-13
c197 1481 0 1.15e-13
c198 1480 0 2.2e-13
c199 1468 0 2.69e-13
c200 77 0 3.13e-13
c201 1465 0 2.76e-13
c202 79 0 4.48e-13
c203 1461 0 4e-11
c204 1460 0 1.1e-13
c205 1459 0 1.15e-13
c206 1458 0 2.2e-13
c207 697 0 5.29e-13
c208 731 0 5.15e-13
c209 734 0 5.37e-13
c210 768 0 5.21e-13
c211 771 0 5.43e-13
c212 805 0 5.31e-13
c213 808 0 5.53e-13
c214 1331 0 3.67e-13
c215 1329 0 2.33e-13
c216 319 0 2.66e-13
c217 1252 0 1.01e-13
c218 315 0 2.6e-13
c219 1243 0 1.15e-13
c220 311 0 2.52e-13
c221 1234 0 1.2e-13
c222 1065 0 1.09e-13
c223 1025 0 1.3e-13
c224 1064 0 1.09e-13
c225 1024 0 1.22e-13
c226 1081 0 1.04e-13
c227 1041 0 1.25e-13
c228 1160 0 1.02e-13
c229 1080 0 1.03e-13
c230 1040 0 1.15e-13
c231 1090 0 1.04e-13
c232 1050 0 1.24e-13
c233 1089 0 1.13e-13
c234 1049 0 1.32e-13
c235 295 0 2.67e-13
c236 299 0 3.03e-13
c237 303 0 3.33e-13
c238 1153 0 1.66e-13
c239 307 0 3.63e-13
c240 1113 0 1.37e-13
c241 1073 0 1.12e-13
c242 290 0 2.56e-13
c243 285 0 2.84e-13
c244 280 0 2.97e-13
c245 873 0 1.62e-13
c246 274 0 3.18e-13
c247 913 0 1.32e-13
c248 953 0 1.08e-13
c249 865 0 1.53e-13
c250 945 0 1.03e-13
c251 905 0 1.26e-13
c252 864 0 1.61e-13
c253 904 0 1.34e-13
c254 944 0 1.06e-13
c255 881 0 1.46e-13
c256 921 0 1.2e-13
c257 880 0 1.53e-13
c258 920 0 1.27e-13
c259 890 0 1.49e-13
c260 970 0 1.01e-13
c261 930 0 1.23e-13
c262 889 0 1.58e-13
c263 929 0 1.32e-13
c264 969 0 1.04e-13
c265 851 0 4.38e-13
c266 852 0 2.03e-13
c267 850 0 1.23e-13
c268 287 0 1.47e-13
c269 849 0 1.21e-13
c270 848 0 1.91e-13
c271 846 0 4e-11
c272 847 0 3.85e-13
c273 844 0 4.38e-13
c274 845 0 2.03e-13
c275 843 0 1.23e-13
c276 292 0 1.32e-13
c277 842 0 1.21e-13
c278 841 0 1.91e-13
c279 839 0 4e-11
c280 840 0 3.85e-13
c281 838 0 4e-11
c282 837 0 1.1e-13
c283 836 0 1.15e-13
c284 835 0 2.2e-13
c285 834 0 4e-11
c286 833 0 1.1e-13
c287 832 0 1.15e-13
c288 831 0 2.2e-13
c289 509 0 1.02e-13
c290 436 0 1.66e-13
c291 433 0 1.37e-13
c292 500 0 1.04e-13
c293 492 0 1.13e-13
c294 516 0 1.04e-13
c295 505 0 1.03e-13
c296 431 0 1.12e-13
c297 533 0 1.09e-13
c298 522 0 1.09e-13
c299 495 0 1.24e-13
c300 490 0 1.32e-13
c301 515 0 1.25e-13
c302 503 0 1.15e-13
c303 532 0 1.3e-13
c304 520 0 1.22e-13
c305 374 0 1.01e-13
c306 361 0 1.04e-13
c307 416 0 1.08e-13
c308 412 0 1.03e-13
c309 399 0 1.06e-13
c310 370 0 1.23e-13
c311 363 0 1.32e-13
c312 389 0 1.2e-13
c313 382 0 1.27e-13
c314 418 0 1.32e-13
c315 408 0 1.26e-13
c316 401 0 1.34e-13
c317 223 0 5.48e-13
c318 209 0 5.57e-13
c319 204 0 5.45e-13
c320 190 0 5.54e-13
c321 185 0 5.46e-13
c322 171 0 5.5e-13
c323 166 0 5.4e-13
c324 151 0 5.49e-13
c325 146 0 5.32e-13
c326 131 0 5.46e-13
c327 126 0 5.32e-13
c328 111 0 5.4e-13
c329 106 0 5.34e-13
c330 91 0 5.51e-13
c331 86 0 5.41e-13
c332 546 0 5.25e-13
c333 549 0 5.43e-13
c334 583 0 5.22e-13
c335 586 0 5.37e-13
c336 620 0 5.09e-13
c337 623 0 5.28e-13
c338 657 0 5.04e-13
c339 660 0 5.18e-13
c340 694 0 5.07e-13
c341 375 0 1.49e-13
c342 365 0 1.58e-13
c343 394 0 1.46e-13
c344 384 0 1.53e-13
c345 228 0 5.58e-13
c346 421 0 1.62e-13
c347 413 0 1.53e-13
c348 403 0 1.61e-13
c349 28 0 6.57e-13
c350 339 0 1.01e-13
c351 333 0 1.15e-13
c352 325 0 1.23e-13
c353 24 0 3.18e-13
c354 16 0 3.24e-13
c355 8 0 2e-13
c356 317 0 2.37e-13
c357 62 0 1.66e-13
c358 313 0 2.37e-13
c359 70 0 1.52e-13
c360 309 0 2.34e-13
c361 243 0 1.37e-13
c362 305 0 3.51e-13
c363 251 0 1.22e-13
c364 301 0 3.3e-13
c365 259 0 1.07e-13
c366 297 0 3.04e-13
c367 293 0 2.76e-13
c368 288 0 2.72e-13
c369 283 0 3.06e-13
c370 278 0 3.26e-13
c371 271 0 3.57e-13
c372 275 0 1.65e-13
c373 273 0 2.31e-13
c374 269 0 4.38e-13
c375 270 0 2.03e-13
c376 268 0 1.23e-13
c377 267 0 1.18e-13
c378 266 0 1.21e-13
c379 265 0 1.91e-13
c380 263 0 4e-11
c381 264 0 3.85e-13
c382 261 0 4.38e-13
c383 262 0 2.03e-13
c384 260 0 1.23e-13
c385 258 0 1.21e-13
c386 257 0 1.91e-13
c387 255 0 4e-11
c388 256 0 3.85e-13
c389 253 0 4.38e-13
c390 254 0 2.03e-13
c391 252 0 1.23e-13
c392 250 0 1.21e-13
c393 249 0 1.91e-13
c394 247 0 4e-11
c395 248 0 3.85e-13
c396 245 0 4.38e-13
c397 246 0 2.03e-13
c398 244 0 1.23e-13
c399 242 0 1.21e-13
c400 241 0 1.91e-13
c401 239 0 4e-11
c402 240 0 3.85e-13
c403 238 0 4e-11
c404 237 0 1.1e-13
c405 236 0 1.15e-13
c406 235 0 2.2e-13
c407 34 0 2.83e-13
c408 72 0 4.38e-13
c409 73 0 2.03e-13
c410 71 0 1.23e-13
c411 69 0 1.21e-13
c412 68 0 1.91e-13
c413 66 0 4e-11
c414 67 0 3.85e-13
c415 64 0 4.38e-13
c416 65 0 2.03e-13
c417 63 0 1.23e-13
c418 61 0 1.21e-13
c419 60 0 1.91e-13
c420 58 0 4e-11
c421 59 0 3.85e-13
c422 57 0 4e-11
c423 56 0 1.1e-13
c424 55 0 1.15e-13
c425 54 0 2.2e-13
c426 52 0 4e-11
c427 51 0 1.1e-13
c428 50 0 1.15e-13
c429 49 0 2.2e-13
c430 47 0 4e-11
c431 46 0 1.1e-13
c432 45 0 1.15e-13
c433 44 0 2.2e-13
c434 42 0 4e-11
c435 41 0 1.1e-13
c436 40 0 1.15e-13
c437 39 0 2.2e-13
c438 37 0 4e-11
c439 36 0 1.1e-13
c440 33 0 2.12e-13
c441 35 0 1.15e-13
c442 32 0 4e-11
c443 31 0 1.1e-13
c444 30 0 1.15e-13
c445 29 0 2.2e-13
c446 26 0 4.38e-13
c447 27 0 2.03e-13
c448 25 0 1.23e-13
c449 23 0 1.21e-13
c450 22 0 1.91e-13
c451 20 0 4e-11
c452 21 0 3.85e-13
c453 18 0 4.38e-13
c454 19 0 2.03e-13
c455 17 0 1.23e-13
c456 15 0 1.21e-13
c457 14 0 1.91e-13
c458 12 0 4e-11
c459 13 0 3.85e-13
c460 10 0 4.38e-13
c461 11 0 2.03e-13
c462 9 0 1.23e-13
c463 7 0 1.21e-13
c464 6 0 1.91e-13
c465 4 0 4e-11
c466 5 0 3.85e-13
rin 1 3 0.001
VPHI 1686 0 pwl (0 5 2.5e-08 5 2.6e-08 0 5e-08 0  5.1e-08 5 7.5e-08 5 7.6e-08 0 1e-07 0  1.01e-07 5 1.25e-07 5 1.26e-07 0 1.5e-07 0  1.51e-07 5 1.75e-07 5 1.76e-07 0 2e-07 0  2.01e-07 5 2.25e-07 5 2.26e-07 0 2.5e-07 0  2.51e-07 5 2.75e-07 5 2.76e-07 0 3e-07 0  3.01e-07 5 3.25e-07 5 3.26e-07 0 3.5e-07 0  3.51e-07 5 3.75e-07 5 3.76e-07 0 4e-07 0  4.01e-07 5 4.25e-07 5 4.26e-07 0 4.5e-07 0  4.51e-07 5 4.75e-07 5 4.76e-07 0 5e-07 0  5.01e-07 5 )
VMRST 37 0 pwl (0 5 5e-08 5 1e-07 5 1.5e-07 5  2e-07 5 2.5e-07 5 3e-07 5 3.5e-07 5  4e-07 5 4.5e-07 5 5e-07 5 )
VENVOTER#1 32 0 pwl (0 5 5e-08 5 1e-07 5 1.5e-07 5  2e-07 5 2.5e-07 5 3e-07 5 3.5e-07 5  4e-07 5 4.5e-07 5 5e-07 5 )
VENVOTER#2 1675 0 pwl (0 5 5e-08 5 1e-07 5 1.5e-07 5  2e-07 5 2.5e-07 5 3e-07 5 3.5e-07 5  4e-07 5 4.5e-07 5 5e-07 5 )
VBSEL#0 1483 0 pwl (0 0 5e-08 0 5.1e-08 5 1e-07 5  1.01e-07 0 1.5e-07 0 1.51e-07 5 2.5e-07 5  2.51e-07 0 3e-07 0 3.01e-07 5 4.5e-07 5  4.51e-07 0 5e-07 0 5.01e-07 5 )
VBSEL#1 1487 0 pwl (0 0 1e-07 0 1.01e-07 5 2e-07 5  2.01e-07 0 2.5e-07 0 2.51e-07 5 3.5e-07 5  3.51e-07 0 4e-07 0 4.01e-07 5 4.5e-07 5  4.51e-07 0 5.5e-07 0 )
VIN#7 1461 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#6 838 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#5 834 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#4 238 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#3 57 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#2 52 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#1 47 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VIN#0 42 0 pwl (0 5 2e-07 5 2.01e-07 0 3.5e-07 0  3.51e-07 5 4.5e-07 5 6.5e-07 5 )
VINBAR#7 1491 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#6 1495 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#5 1660 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#4 1664 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#3 1709 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#2 1705 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#1 1701 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VINBAR#0 1697 0 pwl (0 0 2e-07 0 2.01e-07 5 3.5e-07 5  3.51e-07 0 4.5e-07 0 6.5e-07 0 )
VVDD 1 0 5
.temp 125 
*.print TRAN v(1686) v(1665) v(1496) v(846) v(839) v(263) v(255) v(247) v(239) v(66) v(58) v(4) 
.options limpts=50000 itl5=50000
*.TRAN 1e-09 5e-07
.op
.end
