REGULATOR  2001.05.26 Y.INOUE
*.OP
*.OPTIONS NOMOD
*.OPTIONS CONV=4:#ITER=361 CONV=1:#ITER=153 CONV=2:#ITER=127 CONV=3:NOCON
*.OPTIONS CONV=2 
VCC 1 0 DC 5.0
*VCC 1 0 DC 3.5
RLOAD 22 0 420.0
R1 2 22 29.6K
R2 2 0 12.0K
R3 1 3 10.0K
R4 6 22 2.0K
R5 7 0 30.0K
R6 10 0 10.0K
R7 11 22 11.0K
R8 11 14 10.0K
R9 13 0 560.0
R10 9 11 10.0K
R11 15 22 15.0K
R12 15 0 10.0K
R13 16 18 10.0K
R14 20 0 5.0K
R15 1 21 100K
Q1 22 3 1 QP 28
Q2 0 4 3 QP 3
Q3 1 8 4 QN
Q4 4 9 0 QN
Q5 5 2 7 QN 2
Q6 8 11 7 QN 2
Q7 5 5 1 QP
Q8 8 5 1 QP
Q9 22 6 8 QP
Q10 10 10 11 QP
Q11 12 10 11 QP
Q12 12 14 0 QN
Q13 0 12 11 QP
Q14 14 9 13 QN 3
Q15 9 9 0 QN
Q16 4 17 0 QN
Q17 17 17 0 QN
Q18 16 16 17 QN
Q19 1 15 20 QN
Q20 19 16 20 QN
Q21 19 21 20 QN
Q22 18 19 1 QP
Q23 19 19 1 QP
Q24 21 21 0 QN
.MODEL QN NPN (IS=1.0E-16 BF=80 BR=1 VA=50 RE=10 RB=100 RC=1K)
.MODEL QP PNP (IS=1.0E-15 BF=80 BR=1 VA=50 RE=10 RB=100 RC=10)
*.END

.OPTIONS DELMAX=1000ns
.op
*.pstran convval=1.0e-05 initstep=1.0e-05 minstep=1.0e-09 maxstep=1.0e+6 tau=1.0e-05 vbe0=0.0 kvgs0=0.0  tauramp=0.0
.end