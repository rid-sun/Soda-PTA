MOSMEM - MOS MEMORY CELL
.WIDTH IN=72
*.OPT ABSTOL=1U
*.OPT ACCT LIST NODE
*.TRAN 20NS 2US
VDD 9 0 DC 5
VS 7 0 PULSE(2 0 520NS 20NS 20NS 500NS 2000NS)
VW 1 0 PULSE(0 2 20NS 20NS 500NS 200NS)
VWB 2 0 PULSE(2 0 20NS 20NS 20NS 2000NS 2000NS)
M1 3 1 0 0 MOD W=250U L=5U
M2 4 2 0 0 MOD W=250U L=5U
M3 9 9 3 0 MOD W=5U   L=5U
M4 9 9 4 0 MOD W=5U   L=5U
M5 5 7 3 0 MOD W=50U  L=5U
M6 6 7 4 0 MOD W=50U  L=5U
M7 5 6 0 0 MOD W=250U  L=5U
M8 6 5 0 0 MOD W=250U  L=5U
M9 9 9 5 0 MOD W=5U   L=5U
M10 9 9 6 0 MOD W=5U  L=5U
M11 8 4 0 0 MOD W=250U L=5U
M12 9 9 8 0 MOD W=5U   L=5U
.MODEL MOD NMOS(VTO=0.5 PHI=0.7 KP=1.0E-6 GAMMA=1.83 LAMBDA=0.115
+   LEVEL=1 CGSO=1U CGDO=1U CBD=50P CBS=50P)
*.PRINT DC V(5) V(6)
*.PLOT DC V(6)
*.PLOT TRAN V(6) V(5) V(7) V(1) V(2)
*.END


.OPTIONS DELMAX=1000ns
.op
*.pstran convval=1.0e-05 initstep=1.0e-05 minstep=1.0e-06 maxstep=1.0e6 tau=1.0e-04 vbe0=0.0 kvgs0=0.0  tauramp=0.0
.end 