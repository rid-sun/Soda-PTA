DIFFICULT CIRCUIT Y.I 2001.5.28
*.OP
*.OPTIONS NOMOD
VCC 1 0 DC 3.3
R1 1 4 50
R2 4 0 50
R3 1 2 20
R4 1 3 1
R5 6 7 20
R6 7 0 100
R7 4 8 200
R8 4 9 200
Q1 2 4 5 QN 
Q2 3 4 5 QN 
Q3 5 5 0 QN 
Q4 6 2 1 QP 
Q5 8 7 0 QN 
Q6 9 3 1 QP 
.MODEL QN NPN (IS=1.0E-14 BF=100
.MODEL QP PNP (IS=1.0E-14 BF=100
*.END
.OPTIONS DELMAX=1000ns
.op
*.gmin
.end