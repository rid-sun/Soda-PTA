add32.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.62249   kp = 6.32664e-05   gamma = 0.639243
+   phi = 0.31
+
+   cgso = 2.89e-10   cgdo = 2.89e-10
+   rsh = 60   cj = 0.000327
+   mj = 1.067   cjsw = 1.74e-10   mjsw = 0.195
+   tox = 2.25e-08   nsub = 1.066e+16
+   nss = 3e+10   nfs = 4.55168e+12   tpg = 1
+   xj = 9e-07   ld = 0   uo = 1215.74
+   ucrit = 174667   uexp = 0.0461235
+   vmax = 177269   neff = 4.6883
+
+   delta = 0
.model penh pmos
+ level = 2
+   vto = -0.63025   kp = 2.63544e-05   gamma = 0.618101
+   phi = 0.541111
+
+   cgso = 3.35e-10   cgdo = 3.35e-10
+   rsh = 150   cj = 0.000475
+   mj = 0.341   cjsw = 2.23e-10   mjsw = 0.307
+   tox = 2.25e-08   nsub = 6.57544e+16
+   nss = 3e+10   nfs = 1.66844e+11   tpg = -1
+   xj = 1.12799e-07   ld = 3e-08   uo = 361.941
+   ucrit = 637449   uexp = 0.0888696
+   vmax = 63253.3   neff = 0.64354
+
+   delta = 0
.subckt add 1 2 3 4 5
+ 6 7
m1 7 8 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m2 7 8 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m3 9 10 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd20 8 10 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m4 2 11 8 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m5 8 11 9 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m6 11 12 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m7 12 3 13 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m8 13 4 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m9 11 12 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd9 1 3 12 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m10 12 4 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m11 10 14 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd7 1 5 14 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m12 14 15 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m13 10 14 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m14 16 15 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m15 6 17 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m16 6 17 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m17 18 19 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd5 17 19 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m18 2 20 17 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd6 17 20 18 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m19 21 5 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m20 19 22 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd3 1 15 22 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m21 22 21 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m22 19 22 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m23 22 15 23 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m24 23 21 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m25 21 5 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m26 24 15 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m27 20 25 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd4 1 5 25 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m28 25 24 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m29 20 25 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m30 25 5 26 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m31 26 24 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m32 24 15 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m33 27 4 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd1 1 3 28 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m34 28 27 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m35 29 28 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m36 28 3 30 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
m37 27 4 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd28 15 31 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd27 15 31 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd26 32 29 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd25 31 29 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd23 2 33 31 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd19 31 33 32 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd18 33 34 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd17 34 4 35 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd16 35 36 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd15 36 3 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd14 33 34 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd13 1 4 34 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd12 34 36 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd11 36 3 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd8 29 28 1 1 penh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd2 30 27 2 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
mXd10 14 5 16 2 nenh l=8e-07 w=3.2e-06 
+ as=1.28e-11 ad=1.28e-11 ps=1.44e-05 pd=1.44e-05 
csum 6 2 3.46e-15
cb 4 2 2.611e-14
ca 3 2 2.534e-14
ccout 7 2 4.99e-15
cc 5 2 2.304e-14
cI0 8 2 3.84e-15
cI2 11 2 3.46e-15
cI3 12 2 3.84e-15
cI5 10 2 4.99e-15
cI6 14 2 4.61e-15
cI8 28 2 3.84e-15
cI9 17 2 3.84e-15
cI11 19 2 5.38e-15
cI12 22 2 4.61e-15
cI13 15 2 1.114e-14
cI14 21 2 5.38e-15
cI16 20 2 5.57e-15
cI17 25 2 4.61e-15
cI18 24 2 6.14e-15
cI20 27 2 5.38e-15
cI22 31 2 3.84e-15
cI23 29 2 5.38e-15
cI25 33 2 3.46e-15
cI26 34 2 3.84e-15
cI28 36 2 3.07e-15
.ends add
xaddX1 1 0 3 4 5
+ 6 7 add
xaddX2 1 0 37 38 7
+ 39 40 add
xaddX3 1 0 70 71 40
+ 72 73 add
xaddX4 1 0 103 104 73
+ 105 106 add
xaddX5 1 0 136 137 106
+ 138 139 add
xaddX6 1 0 169 170 139
+ 171 172 add
xaddX7 1 0 202 203 172
+ 204 205 add
xaddX8 1 0 235 236 205
+ 237 238 add
xaddX9 1 0 268 269 238
+ 270 271 add
xaddX10 1 0 301 302 271
+ 303 304 add
xaddX11 1 0 334 335 304
+ 336 337 add
xaddX12 1 0 367 368 337
+ 369 370 add
xaddX13 1 0 400 401 370
+ 402 403 add
xaddX14 1 0 433 434 403
+ 435 436 add
xaddX15 1 0 466 467 436
+ 468 469 add
xaddX16 1 0 499 500 469
+ 501 502 add
xaddY1 1 0 532 533 502
+ 534 535 add
xaddY2 1 0 565 566 535
+ 567 568 add
xaddY3 1 0 598 599 568
+ 600 601 add
xaddY4 1 0 631 632 601
+ 633 634 add
xaddY5 1 0 664 665 634
+ 666 667 add
xaddY6 1 0 697 698 667
+ 699 700 add
xaddY7 1 0 730 731 700
+ 732 733 add
xaddY8 1 0 763 764 733
+ 765 766 add
xaddY9 1 0 796 797 766
+ 798 799 add
xaddY10 1 0 829 830 799
+ 831 832 add
xaddY11 1 0 862 863 832
+ 864 865 add
xaddY12 1 0 895 896 865
+ 897 898 add
xaddY13 1 0 928 929 898
+ 930 931 add
xaddY14 1 0 961 962 931
+ 963 964 add
xaddY15 1 0 994 995 964
+ 996 997 add
xaddY16 1 0 1027 1028 997
+ 1029 1030 add
Va1 3 0 pwl (0 0 2e-08 0 2.1e-08 5 4e-08 5 
+ 4.1e-08 0 5e-08 0 5.1e-08 5 7e-08 5 
+ 7.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.7e-07 0 1.71e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.9e-07 0 2.91e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.8e-07 0 3.81e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.2e-07 0 4.21e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 4.7e-07 5 
+ 4.71e-07 0 5.3e-07 0 5.31e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6e-07 0 6.01e-07 5 6.4e-07 5 
+ 6.41e-07 0 6.9e-07 0 6.91e-07 5 7e-07 5 
+ 7.01e-07 0 7.3e-07 0 7.31e-07 5 7.5e-07 5 
+ 7.51e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.9e-07 0 8.91e-07 5 9e-07 5 
+ 9.01e-07 0 9.2e-07 0 9.21e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.6e-07 0 9.61e-07 5 9.8e-07 5 
+ 9.81e-07 0 1e-06 0 )
Va2 37 0 pwl (0 5 1e-08 5 1.1e-08 0 4e-08 0 
+ 4.1e-08 5 5e-08 5 5.1e-08 0 7e-08 0 
+ 7.1e-08 5 9e-08 5 9.1e-08 0 1.1e-07 0 
+ 1.11e-07 5 1.2e-07 5 1.21e-07 0 1.3e-07 0 
+ 1.31e-07 5 1.4e-07 5 1.41e-07 0 1.7e-07 0 
+ 1.71e-07 5 2.3e-07 5 2.31e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.5e-07 5 2.51e-07 0 2.7e-07 0 
+ 2.71e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.3e-07 5 3.31e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.9e-07 5 3.91e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.5e-07 5 4.51e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.9e-07 5 4.91e-07 0 5e-07 0 
+ 5.01e-07 5 5.2e-07 5 5.21e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.9e-07 5 5.91e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.3e-07 5 6.31e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.8e-07 5 6.81e-07 0 7e-07 0 
+ 7.01e-07 5 7.1e-07 5 7.11e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.6e-07 5 7.61e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.8e-07 5 7.81e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.4e-07 5 8.41e-07 0 8.6e-07 0 
+ 8.61e-07 5 8.7e-07 5 8.71e-07 0 8.9e-07 0 
+ 8.91e-07 5 9e-07 5 9.01e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.2e-07 5 9.21e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 1e-06 5 1.01e-06 5 )
Va3 70 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 5e-08 5 5.1e-08 0 8e-08 0 
+ 8.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 2e-07 0 
+ 2.01e-07 5 2.1e-07 5 2.11e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.9e-07 5 2.91e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.3e-07 5 3.31e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.9e-07 5 3.91e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.3e-07 5 4.31e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.5e-07 5 4.51e-07 0 4.7e-07 0 
+ 4.71e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.4e-07 5 5.41e-07 0 5.5e-07 0 
+ 5.51e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.8e-07 5 5.81e-07 0 6e-07 0 
+ 6.01e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.4e-07 5 6.41e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.7e-07 5 6.71e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.5e-07 5 7.51e-07 0 7.9e-07 0 
+ 7.91e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.6e-07 5 8.61e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.02e-06 5 )
Va4 103 0 pwl (0 0 2e-08 0 2.1e-08 5 5e-08 5 
+ 5.1e-08 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.3e-07 0 1.31e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.7e-07 5 
+ 1.71e-07 0 1.8e-07 0 1.81e-07 5 2e-07 5 
+ 2.01e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.6e-07 0 2.61e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 4e-07 5 
+ 4.01e-07 0 4.1e-07 0 4.11e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.5e-07 0 4.51e-07 5 4.7e-07 5 
+ 4.71e-07 0 4.9e-07 0 4.91e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.8e-07 0 5.81e-07 5 6e-07 5 
+ 6.01e-07 0 6.1e-07 0 6.11e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.7e-07 0 6.71e-07 5 6.9e-07 5 
+ 6.91e-07 0 7.1e-07 0 7.11e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.3e-07 0 7.31e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.9e-07 0 7.91e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.9e-07 0 8.91e-07 5 9e-07 5 
+ 9.01e-07 0 9.1e-07 0 9.11e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 1e-06 0 1.02e-06 0 )
Va5 136 0 pwl (0 5 1e-08 5 1.1e-08 0 3e-08 0 
+ 3.1e-08 5 6e-08 5 6.1e-08 0 7e-08 0 
+ 7.1e-08 5 9e-08 5 9.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.8e-07 5 1.81e-07 0 1.9e-07 0 
+ 1.91e-07 5 2e-07 5 2.01e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.8e-07 5 2.81e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.9e-07 5 3.91e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.2e-07 5 4.21e-07 0 4.8e-07 0 
+ 4.81e-07 5 5.1e-07 5 5.11e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.4e-07 5 5.41e-07 0 5.5e-07 0 
+ 5.51e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.3e-07 5 6.31e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.7e-07 5 6.71e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.2e-07 5 7.21e-07 0 7.3e-07 0 
+ 7.31e-07 5 7.4e-07 5 7.41e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.7e-07 5 7.71e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.7e-07 5 8.71e-07 0 8.9e-07 0 
+ 8.91e-07 5 9e-07 5 9.01e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.2e-07 5 9.21e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.4e-07 5 9.41e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.6e-07 5 9.61e-07 0 1e-06 0 
+ 1.001e-06 5 1.01e-06 5 )
Va6 169 0 pwl (0 5 3e-08 5 3.1e-08 0 5e-08 0 
+ 5.1e-08 5 8e-08 5 8.1e-08 0 1.3e-07 0 
+ 1.31e-07 5 1.4e-07 5 1.41e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.8e-07 5 1.81e-07 0 1.9e-07 0 
+ 1.91e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.3e-07 5 2.31e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.7e-07 5 2.71e-07 0 3e-07 0 
+ 3.01e-07 5 3.4e-07 5 3.41e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 3.8e-07 0 
+ 3.81e-07 5 3.9e-07 5 3.91e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.3e-07 5 4.31e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.7e-07 5 4.71e-07 0 4.8e-07 0 
+ 4.81e-07 5 5e-07 5 5.01e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.9e-07 5 5.91e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.6e-07 5 6.61e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.8e-07 5 6.81e-07 0 7e-07 0 
+ 7.01e-07 5 7.2e-07 5 7.21e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.6e-07 5 7.61e-07 0 7.7e-07 0 
+ 7.71e-07 5 8.4e-07 5 8.41e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.9e-07 5 8.91e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.2e-07 5 9.21e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.6e-07 5 9.61e-07 0 9.8e-07 0 
+ 9.81e-07 5 1e-06 5 1.03e-06 5 )
Va7 202 0 pwl (0 5 3e-08 5 3.1e-08 0 4e-08 0 
+ 4.1e-08 5 6e-08 5 6.1e-08 0 7e-08 0 
+ 7.1e-08 5 8e-08 5 8.1e-08 0 9e-08 0 
+ 9.1e-08 5 1e-07 5 1.01e-07 0 1.3e-07 0 
+ 1.31e-07 5 1.4e-07 5 1.41e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 1.9e-07 0 
+ 1.91e-07 5 2.7e-07 5 2.71e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.8e-07 5 3.81e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.2e-07 5 4.21e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.4e-07 5 4.41e-07 0 5e-07 0 
+ 5.01e-07 5 5.1e-07 5 5.11e-07 0 5.2e-07 0 
+ 5.21e-07 5 5.3e-07 5 5.31e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.8e-07 5 5.81e-07 0 5.9e-07 0 
+ 5.91e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.5e-07 5 6.51e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.7e-07 5 6.71e-07 0 6.8e-07 0 
+ 6.81e-07 5 6.9e-07 5 6.91e-07 0 7e-07 0 
+ 7.01e-07 5 7.7e-07 5 7.71e-07 0 7.9e-07 0 
+ 7.91e-07 5 8e-07 5 8.01e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.6e-07 5 8.61e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.6e-07 5 9.61e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Va8 235 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 4e-08 5 4.1e-08 0 1.2e-07 0 
+ 1.21e-07 5 1.4e-07 5 1.41e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.3e-07 5 2.31e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.7e-07 5 2.71e-07 0 3e-07 0 
+ 3.01e-07 5 3.1e-07 5 3.11e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 3.8e-07 0 
+ 3.81e-07 5 4.1e-07 5 4.11e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.4e-07 5 4.41e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.7e-07 5 4.71e-07 0 4.9e-07 0 
+ 4.91e-07 5 5e-07 5 5.01e-07 0 5.2e-07 0 
+ 5.21e-07 5 5.3e-07 5 5.31e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.8e-07 5 5.81e-07 0 5.9e-07 0 
+ 5.91e-07 5 6e-07 5 6.01e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.5e-07 5 6.51e-07 0 6.8e-07 0 
+ 6.81e-07 5 6.9e-07 5 6.91e-07 0 7e-07 0 
+ 7.01e-07 5 7.3e-07 5 7.31e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.8e-07 5 7.81e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 9e-07 5 9.01e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 9.9e-07 0 
+ 9.91e-07 5 1e-06 5 )
Va9 268 0 pwl (0 0 1e-08 0 1.1e-08 5 3e-08 5 
+ 3.1e-08 0 4e-08 0 4.1e-08 5 5e-08 5 
+ 5.1e-08 0 8e-08 0 8.1e-08 5 1.1e-07 5 
+ 1.11e-07 0 1.3e-07 0 1.31e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.6e-07 0 2.61e-07 5 2.7e-07 5 
+ 2.71e-07 0 3e-07 0 3.01e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 3.8e-07 5 
+ 3.81e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.4e-07 0 4.41e-07 5 4.8e-07 5 
+ 4.81e-07 0 5e-07 0 5.01e-07 5 5.1e-07 5 
+ 5.11e-07 0 5.4e-07 0 5.41e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.7e-07 0 5.71e-07 5 5.8e-07 5 
+ 5.81e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.9e-07 0 6.91e-07 5 7e-07 5 
+ 7.01e-07 0 7.1e-07 0 7.11e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 8.3e-07 0 8.31e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.5e-07 0 8.51e-07 5 8.6e-07 5 
+ 8.61e-07 0 8.9e-07 0 8.91e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.4e-07 0 9.41e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.7e-07 0 9.71e-07 5 9.9e-07 5 
+ 9.91e-07 0 1e-06 0 1.01e-06 0 )
Va10 301 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 4e-08 5 
+ 4.1e-08 0 5e-08 0 5.1e-08 5 7e-08 5 
+ 7.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.2e-07 0 1.21e-07 5 1.3e-07 5 
+ 1.31e-07 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 2e-07 0 2.01e-07 5 2.1e-07 5 
+ 2.11e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.7e-07 0 2.71e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.3e-07 0 4.31e-07 5 4.4e-07 5 
+ 4.41e-07 0 4.6e-07 0 4.61e-07 5 4.7e-07 5 
+ 4.71e-07 0 4.9e-07 0 4.91e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.4e-07 0 5.41e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.1e-07 0 6.11e-07 5 6.8e-07 5 
+ 6.81e-07 0 7e-07 0 7.01e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.3e-07 0 7.31e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.8e-07 0 7.81e-07 5 7.9e-07 5 
+ 7.91e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.6e-07 0 8.61e-07 5 8.9e-07 5 
+ 8.91e-07 0 9.1e-07 0 9.11e-07 5 9.6e-07 5 
+ 9.61e-07 0 1e-06 0 1.01e-06 0 )
Va11 334 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 7e-08 5 
+ 7.1e-08 0 8e-08 0 8.1e-08 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.9e-07 0 1.91e-07 5 2e-07 5 
+ 2.01e-07 0 2.1e-07 0 2.11e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.3e-07 0 3.31e-07 5 3.5e-07 5 
+ 3.51e-07 0 4e-07 0 4.01e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.2e-07 0 4.21e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.4e-07 0 4.41e-07 5 4.7e-07 5 
+ 4.71e-07 0 5.1e-07 0 5.11e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.5e-07 0 5.51e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.8e-07 0 5.81e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.7e-07 0 6.71e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.9e-07 5 
+ 7.91e-07 0 8e-07 0 8.01e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.4e-07 0 8.41e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 8.9e-07 5 
+ 8.91e-07 0 9e-07 0 9.01e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.3e-07 0 9.31e-07 5 9.4e-07 5 
+ 9.41e-07 0 9.5e-07 0 9.51e-07 5 9.8e-07 5 
+ 9.81e-07 0 1e-06 0 )
Va12 367 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 5e-08 5 5.1e-08 0 8e-08 0 
+ 8.1e-08 5 1e-07 5 1.01e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.6e-07 5 1.61e-07 0 1.9e-07 0 
+ 1.91e-07 5 2.1e-07 5 2.11e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.7e-07 5 2.71e-07 0 2.8e-07 0 
+ 2.81e-07 5 3.4e-07 5 3.41e-07 0 3.8e-07 0 
+ 3.81e-07 5 4.1e-07 5 4.11e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.2e-07 5 5.21e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.8e-07 0 
+ 5.81e-07 5 5.9e-07 5 5.91e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.3e-07 5 7.31e-07 0 7.6e-07 0 
+ 7.61e-07 5 8e-07 5 8.01e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.9e-07 5 8.91e-07 0 9e-07 0 
+ 9.01e-07 5 9.1e-07 5 9.11e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.5e-07 5 9.51e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 9.9e-07 0 
+ 9.91e-07 5 1e-06 5 )
Va13 400 0 pwl (0 0 3e-08 0 3.1e-08 5 4e-08 5 
+ 4.1e-08 0 5e-08 0 5.1e-08 5 6e-08 5 
+ 6.1e-08 0 7e-08 0 7.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.5e-07 0 1.51e-07 5 1.7e-07 5 
+ 1.71e-07 0 1.8e-07 0 1.81e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.6e-07 0 2.61e-07 5 2.7e-07 5 
+ 2.71e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 4e-07 0 4.01e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.2e-07 0 4.21e-07 5 4.6e-07 5 
+ 4.61e-07 0 4.7e-07 0 4.71e-07 5 4.8e-07 5 
+ 4.81e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.5e-07 0 5.51e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.8e-07 0 6.81e-07 5 7e-07 5 
+ 7.01e-07 0 7.3e-07 0 7.31e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 8.1e-07 0 8.11e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.7e-07 0 8.71e-07 5 8.8e-07 5 
+ 8.81e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 9.5e-07 5 
+ 9.51e-07 0 1e-06 0 1.03e-06 0 )
Va14 433 0 pwl (0 0 1e-08 0 1.1e-08 5 3e-08 5 
+ 3.1e-08 0 4e-08 0 4.1e-08 5 7e-08 5 
+ 7.1e-08 0 1e-07 0 1.01e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 2.1e-07 0 2.11e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.4e-07 0 2.41e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.6e-07 0 2.61e-07 5 2.8e-07 5 
+ 2.81e-07 0 2.9e-07 0 2.91e-07 5 3e-07 5 
+ 3.01e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.8e-07 0 3.81e-07 5 4e-07 5 
+ 4.01e-07 0 4.2e-07 0 4.21e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.5e-07 0 4.51e-07 5 4.7e-07 5 
+ 4.71e-07 0 4.8e-07 0 4.81e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.1e-07 0 5.11e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.7e-07 0 5.71e-07 5 5.8e-07 5 
+ 5.81e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.9e-07 0 6.91e-07 5 7.1e-07 5 
+ 7.11e-07 0 7.3e-07 0 7.31e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.4e-07 0 8.41e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.6e-07 0 8.61e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 1e-06 0 1.01e-06 0 )
Va15 466 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 4e-08 5 
+ 4.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1e-07 0 1.01e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.3e-07 0 1.31e-07 5 1.5e-07 5 
+ 1.51e-07 0 1.7e-07 0 1.71e-07 5 1.8e-07 5 
+ 1.81e-07 0 2.1e-07 0 2.11e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.4e-07 0 2.41e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.8e-07 0 2.81e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.8e-07 0 3.81e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.2e-07 0 4.21e-07 5 4.4e-07 5 
+ 4.41e-07 0 4.7e-07 0 4.71e-07 5 4.8e-07 5 
+ 4.81e-07 0 5e-07 0 5.01e-07 5 5.1e-07 5 
+ 5.11e-07 0 5.2e-07 0 5.21e-07 5 5.5e-07 5 
+ 5.51e-07 0 6e-07 0 6.01e-07 5 6.6e-07 5 
+ 6.61e-07 0 7.2e-07 0 7.21e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.5e-07 0 8.51e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 9e-07 5 
+ 9.01e-07 0 9.1e-07 0 9.11e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.3e-07 0 9.31e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.7e-07 0 9.71e-07 5 1e-06 5 
+ 1.001e-06 0 1.01e-06 0 )
Va16 499 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 6e-08 0 
+ 6.1e-08 5 8e-08 5 8.1e-08 0 1.1e-07 0 
+ 1.11e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 1.8e-07 5 1.81e-07 0 2e-07 0 
+ 2.01e-07 5 2.2e-07 5 2.21e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.5e-07 0 
+ 3.51e-07 5 3.6e-07 5 3.61e-07 0 3.7e-07 0 
+ 3.71e-07 5 4e-07 5 4.01e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.7e-07 5 4.71e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.4e-07 5 5.41e-07 0 5.9e-07 0 
+ 5.91e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.4e-07 5 6.41e-07 0 6.7e-07 0 
+ 6.71e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.4e-07 5 7.41e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.6e-07 5 7.61e-07 0 7.8e-07 0 
+ 7.81e-07 5 7.9e-07 5 7.91e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.4e-07 5 8.41e-07 0 8.5e-07 0 
+ 8.51e-07 5 8.6e-07 5 8.61e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.9e-07 5 8.91e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.4e-07 5 9.41e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.6e-07 5 9.61e-07 0 9.7e-07 0 
+ 9.71e-07 5 1e-06 5 )
Vb1 4 0 pwl (0 5 1e-08 5 1.1e-08 0 3e-08 0 
+ 3.1e-08 5 5e-08 5 5.1e-08 0 6e-08 0 
+ 6.1e-08 5 7e-08 5 7.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.3e-07 0 
+ 1.31e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 1.9e-07 5 1.91e-07 0 2e-07 0 
+ 2.01e-07 5 2.2e-07 5 2.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.5e-07 5 2.51e-07 0 3e-07 0 
+ 3.01e-07 5 3.1e-07 5 3.11e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.6e-07 5 3.61e-07 0 3.8e-07 0 
+ 3.81e-07 5 3.9e-07 5 3.91e-07 0 4e-07 0 
+ 4.01e-07 5 4.2e-07 5 4.21e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.6e-07 5 4.61e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.3e-07 5 5.31e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.6e-07 5 5.61e-07 0 5.8e-07 0 
+ 5.81e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.8e-07 5 6.81e-07 0 6.9e-07 0 
+ 6.91e-07 5 7.1e-07 5 7.11e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.5e-07 5 7.51e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.7e-07 5 7.71e-07 0 7.9e-07 0 
+ 7.91e-07 5 8e-07 5 8.01e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.6e-07 5 8.61e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.8e-07 5 8.81e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.01e-06 5 )
Vb2 38 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 4e-08 0 4.1e-08 5 6e-08 5 
+ 6.1e-08 0 1.1e-07 0 1.11e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.7e-07 0 1.71e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.3e-07 0 2.31e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.5e-07 0 3.51e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.5e-07 0 4.51e-07 5 4.9e-07 5 
+ 4.91e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.4e-07 0 5.41e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.6e-07 0 5.61e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.9e-07 0 6.91e-07 5 7e-07 5 
+ 7.01e-07 0 7.3e-07 0 7.31e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.8e-07 0 7.81e-07 5 7.9e-07 5 
+ 7.91e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.5e-07 0 9.51e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 1.01e-06 0 )
Vb3 71 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 7e-08 0 
+ 7.1e-08 5 9e-08 5 9.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.7e-07 0 
+ 1.71e-07 5 2.2e-07 5 2.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.6e-07 5 2.61e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 3.9e-07 0 
+ 3.91e-07 5 4e-07 5 4.01e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.9e-07 5 4.91e-07 0 5e-07 0 
+ 5.01e-07 5 5.1e-07 5 5.11e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.5e-07 5 5.51e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.8e-07 5 5.81e-07 0 5.9e-07 0 
+ 5.91e-07 5 6.2e-07 5 6.21e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.9e-07 5 6.91e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.5e-07 5 7.51e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.9e-07 5 7.91e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.5e-07 5 8.51e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9e-07 0 
+ 9.01e-07 5 9.1e-07 5 9.11e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.02e-06 5 )
Vb4 104 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 4e-08 5 4.1e-08 0 6e-08 0 
+ 6.1e-08 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.4e-07 5 1.41e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 2.2e-07 5 2.21e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.9e-07 5 3.91e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.3e-07 5 4.31e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.6e-07 5 4.61e-07 0 4.8e-07 0 
+ 4.81e-07 5 5e-07 5 5.01e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 6e-07 0 
+ 6.01e-07 5 6.1e-07 5 6.11e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 7e-07 0 
+ 7.01e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.3e-07 5 7.31e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.5e-07 5 7.51e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.8e-07 5 7.81e-07 0 7.9e-07 0 
+ 7.91e-07 5 8.1e-07 5 8.11e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.8e-07 5 8.81e-07 0 9e-07 0 
+ 9.01e-07 5 9.2e-07 5 9.21e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.7e-07 5 9.71e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vb5 137 0 pwl (0 0 3e-08 0 3.1e-08 5 5e-08 5 
+ 5.1e-08 0 7e-08 0 7.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.5e-07 0 1.51e-07 5 2e-07 5 
+ 2.01e-07 0 2.1e-07 0 2.11e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.8e-07 5 
+ 2.81e-07 0 3e-07 0 3.01e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.5e-07 0 3.51e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 4e-07 5 
+ 4.01e-07 0 4.1e-07 0 4.11e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.4e-07 0 4.41e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.7e-07 0 4.71e-07 5 4.8e-07 5 
+ 4.81e-07 0 5.1e-07 0 5.11e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.6e-07 0 6.61e-07 5 6.7e-07 5 
+ 6.71e-07 0 6.9e-07 0 6.91e-07 5 7.2e-07 5 
+ 7.21e-07 0 8e-07 0 8.01e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.6e-07 0 8.61e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 8.9e-07 5 
+ 8.91e-07 0 9.1e-07 0 9.11e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 1.03e-06 0 )
Vb6 170 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 6e-08 5 6.1e-08 0 7e-08 0 
+ 7.1e-08 5 1e-07 5 1.01e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.6e-07 0 
+ 1.61e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.2e-07 5 2.21e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 3.8e-07 0 
+ 3.81e-07 5 4e-07 5 4.01e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.5e-07 5 4.51e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.7e-07 5 4.71e-07 0 4.8e-07 0 
+ 4.81e-07 5 4.9e-07 5 4.91e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.3e-07 5 5.31e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.8e-07 5 5.81e-07 0 5.9e-07 0 
+ 5.91e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.8e-07 5 6.81e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.2e-07 5 7.21e-07 0 7.3e-07 0 
+ 7.31e-07 5 7.5e-07 5 7.51e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.8e-07 5 7.81e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.4e-07 5 8.41e-07 0 8.8e-07 0 
+ 8.81e-07 5 9e-07 5 9.01e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.2e-07 5 9.21e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.6e-07 0 
+ 9.61e-07 5 1e-06 5 1.02e-06 5 )
Vb7 203 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 6e-08 5 
+ 6.1e-08 0 8e-08 0 8.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.2e-07 0 1.21e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.7e-07 0 1.71e-07 5 1.8e-07 5 
+ 1.81e-07 0 1.9e-07 0 1.91e-07 5 2e-07 5 
+ 2.01e-07 0 2.1e-07 0 2.11e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.4e-07 0 2.41e-07 5 2.7e-07 5 
+ 2.71e-07 0 2.9e-07 0 2.91e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 3.8e-07 5 
+ 3.81e-07 0 4.3e-07 0 4.31e-07 5 4.7e-07 5 
+ 4.71e-07 0 5.2e-07 0 5.21e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.5e-07 0 5.51e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.6e-07 0 6.61e-07 5 6.7e-07 5 
+ 6.71e-07 0 7e-07 0 7.01e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.8e-07 0 7.81e-07 5 7.9e-07 5 
+ 7.91e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.7e-07 0 8.71e-07 5 8.9e-07 5 
+ 8.91e-07 0 9.2e-07 0 9.21e-07 5 9.8e-07 5 
+ 9.81e-07 0 1e-06 0 1.01e-06 0 )
Vb8 236 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 5e-08 5 5.1e-08 0 6e-08 0 
+ 6.1e-08 5 7e-08 5 7.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.2e-07 5 1.21e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.7e-07 5 1.71e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.3e-07 5 2.31e-07 0 2.7e-07 0 
+ 2.71e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.7e-07 0 
+ 3.71e-07 5 3.8e-07 5 3.81e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.5e-07 5 4.51e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.7e-07 5 4.71e-07 0 4.8e-07 0 
+ 4.81e-07 5 4.9e-07 5 4.91e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.4e-07 5 5.41e-07 0 5.5e-07 0 
+ 5.51e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.9e-07 5 5.91e-07 0 6e-07 0 
+ 6.01e-07 5 6.4e-07 5 6.41e-07 0 6.9e-07 0 
+ 6.91e-07 5 7.2e-07 5 7.21e-07 0 7.3e-07 0 
+ 7.31e-07 5 7.5e-07 5 7.51e-07 0 7.8e-07 0 
+ 7.81e-07 5 7.9e-07 5 7.91e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.4e-07 5 8.41e-07 0 8.6e-07 0 
+ 8.61e-07 5 8.7e-07 5 8.71e-07 0 8.9e-07 0 
+ 8.91e-07 5 9.3e-07 5 9.31e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vb9 269 0 pwl (0 0 4e-08 0 4.1e-08 5 1.1e-07 5 
+ 1.11e-07 0 1.3e-07 0 1.31e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.8e-07 5 
+ 1.81e-07 0 1.9e-07 0 1.91e-07 5 2e-07 5 
+ 2.01e-07 0 2.2e-07 0 2.21e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.7e-07 0 2.71e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 4e-07 5 
+ 4.01e-07 0 4.6e-07 0 4.61e-07 5 4.7e-07 5 
+ 4.71e-07 0 4.9e-07 0 4.91e-07 5 5.1e-07 5 
+ 5.11e-07 0 5.2e-07 0 5.21e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.7e-07 0 6.71e-07 5 6.8e-07 5 
+ 6.81e-07 0 6.9e-07 0 6.91e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.6e-07 0 7.61e-07 5 7.9e-07 5 
+ 7.91e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.8e-07 0 8.81e-07 5 9.1e-07 5 
+ 9.11e-07 0 1e-06 0 1.04e-06 0 )
Vb10 302 0 pwl (0 0 1e-08 0 1.1e-08 5 4e-08 5 
+ 4.1e-08 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 1e-07 0 1.01e-07 5 1.1e-07 5 
+ 1.11e-07 0 1.3e-07 0 1.31e-07 5 1.6e-07 5 
+ 1.61e-07 0 2.1e-07 0 2.11e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.4e-07 0 2.41e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.1e-07 0 3.11e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.3e-07 0 4.31e-07 5 4.4e-07 5 
+ 4.41e-07 0 4.5e-07 0 4.51e-07 5 4.7e-07 5 
+ 4.71e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.5e-07 0 5.51e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.2e-07 0 6.21e-07 5 6.5e-07 5 
+ 6.51e-07 0 6.6e-07 0 6.61e-07 5 6.8e-07 5 
+ 6.81e-07 0 8e-07 0 8.01e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.9e-07 0 8.91e-07 5 9.4e-07 5 
+ 9.41e-07 0 9.6e-07 0 9.61e-07 5 9.7e-07 5 
+ 9.71e-07 0 9.8e-07 0 9.81e-07 5 1e-06 5 
+ 1.001e-06 0 1.01e-06 0 )
Vb11 335 0 pwl (0 5 3e-08 5 3.1e-08 0 5e-08 0 
+ 5.1e-08 5 7e-08 5 7.1e-08 0 8e-08 0 
+ 8.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.2e-07 5 1.21e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 2e-07 0 
+ 2.01e-07 5 2.1e-07 5 2.11e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.9e-07 5 2.91e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.2e-07 5 3.21e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.9e-07 0 
+ 3.91e-07 5 4e-07 5 4.01e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.4e-07 5 4.41e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.1e-07 5 5.11e-07 0 5.5e-07 0 
+ 5.51e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 7.4e-07 5 7.41e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.9e-07 5 7.91e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.6e-07 5 8.61e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.8e-07 5 8.81e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.4e-07 5 9.41e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 9.9e-07 0 
+ 9.91e-07 5 1e-06 5 1.03e-06 5 )
Vb12 368 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 8e-08 5 8.1e-08 0 9e-08 0 
+ 9.1e-08 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 1.9e-07 0 
+ 1.91e-07 5 2.1e-07 5 2.11e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.1e-07 5 3.11e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.6e-07 0 
+ 3.61e-07 5 4.4e-07 5 4.41e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.6e-07 5 4.61e-07 0 5e-07 0 
+ 5.01e-07 5 5.3e-07 5 5.31e-07 0 5.4e-07 0 
+ 5.41e-07 5 6.1e-07 5 6.11e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.4e-07 5 6.41e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.7e-07 5 6.71e-07 0 6.9e-07 0 
+ 6.91e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.3e-07 5 7.31e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.6e-07 5 7.61e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.4e-07 5 8.41e-07 0 8.5e-07 0 
+ 8.51e-07 5 8.9e-07 5 8.91e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.2e-07 5 9.21e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.6e-07 5 9.61e-07 0 9.9e-07 0 
+ 9.91e-07 5 1e-06 5 )
Vb13 401 0 pwl (0 0 7e-08 0 7.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.3e-07 0 1.31e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.6e-07 5 
+ 1.61e-07 0 2.2e-07 0 2.21e-07 5 2.6e-07 5 
+ 2.61e-07 0 3.1e-07 0 3.11e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.5e-07 0 3.51e-07 5 3.7e-07 5 
+ 3.71e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.3e-07 0 4.31e-07 5 4.6e-07 5 
+ 4.61e-07 0 5e-07 0 5.01e-07 5 5.1e-07 5 
+ 5.11e-07 0 5.2e-07 0 5.21e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6.1e-07 0 6.11e-07 5 6.8e-07 5 
+ 6.81e-07 0 7.2e-07 0 7.21e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.7e-07 0 7.71e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.6e-07 5 
+ 8.61e-07 0 8.9e-07 0 8.91e-07 5 9e-07 5 
+ 9.01e-07 0 9.1e-07 0 9.11e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 )
Vb14 434 0 pwl (0 0 2e-08 0 2.1e-08 5 4e-08 5 
+ 4.1e-08 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1.3e-07 5 
+ 1.31e-07 0 1.5e-07 0 1.51e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.7e-07 0 1.71e-07 5 1.8e-07 5 
+ 1.81e-07 0 2e-07 0 2.01e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.9e-07 0 2.91e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.7e-07 5 
+ 3.71e-07 0 4e-07 0 4.01e-07 5 4.4e-07 5 
+ 4.41e-07 0 4.5e-07 0 4.51e-07 5 4.6e-07 5 
+ 4.61e-07 0 4.8e-07 0 4.81e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.4e-07 0 5.41e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6.1e-07 0 6.11e-07 5 6.2e-07 5 
+ 6.21e-07 0 6.4e-07 0 6.41e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.8e-07 0 6.81e-07 5 6.9e-07 5 
+ 6.91e-07 0 7.1e-07 0 7.11e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.6e-07 0 8.61e-07 5 8.8e-07 5 
+ 8.81e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.2e-07 0 9.21e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.8e-07 0 9.81e-07 5 9.9e-07 5 
+ 9.91e-07 0 1e-06 0 1.02e-06 0 )
Vb15 467 0 pwl (0 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 7e-08 5 7.1e-08 0 1.1e-07 0 
+ 1.11e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 2e-07 0 
+ 2.01e-07 5 2.1e-07 5 2.11e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.5e-07 5 2.51e-07 0 2.6e-07 0 
+ 2.61e-07 5 3e-07 5 3.01e-07 0 3.5e-07 0 
+ 3.51e-07 5 3.7e-07 5 3.71e-07 0 4e-07 0 
+ 4.01e-07 5 4.1e-07 5 4.11e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.3e-07 5 4.31e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.5e-07 5 4.51e-07 0 4.7e-07 0 
+ 4.71e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5e-07 5 5.01e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.5e-07 5 5.51e-07 0 5.8e-07 0 
+ 5.81e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.5e-07 5 6.51e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.7e-07 5 6.71e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.7e-07 5 7.71e-07 0 7.8e-07 0 
+ 7.81e-07 5 8e-07 5 8.01e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.5e-07 5 8.51e-07 0 8.6e-07 0 
+ 8.61e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 9e-07 5 9.01e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.3e-07 5 9.31e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.7e-07 0 
+ 9.71e-07 5 1e-06 5 1.04e-06 5 )
Vb16 500 0 pwl (0 0 1e-08 0 1.1e-08 5 3e-08 5 
+ 3.1e-08 0 4e-08 0 4.1e-08 5 6e-08 5 
+ 6.1e-08 0 1e-07 0 1.01e-07 5 1.1e-07 5 
+ 1.11e-07 0 1.2e-07 0 1.21e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.9e-07 0 1.91e-07 5 2e-07 5 
+ 2.01e-07 0 2.2e-07 0 2.21e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.5e-07 0 2.51e-07 5 2.7e-07 5 
+ 2.71e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.1e-07 0 3.11e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.3e-07 0 3.31e-07 5 3.4e-07 5 
+ 3.41e-07 0 3.6e-07 0 3.61e-07 5 3.8e-07 5 
+ 3.81e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.4e-07 0 4.41e-07 5 4.7e-07 5 
+ 4.71e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.6e-07 0 6.61e-07 5 6.8e-07 5 
+ 6.81e-07 0 6.9e-07 0 6.91e-07 5 7.1e-07 5 
+ 7.11e-07 0 7.4e-07 0 7.41e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.7e-07 0 7.71e-07 5 8e-07 5 
+ 8.01e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.6e-07 0 8.61e-07 5 8.8e-07 5 
+ 8.81e-07 0 9.2e-07 0 9.21e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.8e-07 0 9.81e-07 5 9.9e-07 5 
+ 9.91e-07 0 1e-06 0 )
Vaa1 532 0 pwl (0 5 5e-08 5 5.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.7e-07 5 1.71e-07 0 1.8e-07 0 
+ 1.81e-07 5 2.1e-07 5 2.11e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.6e-07 5 2.61e-07 0 2.7e-07 0 
+ 2.71e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.2e-07 5 3.21e-07 0 3.7e-07 0 
+ 3.71e-07 5 3.8e-07 5 3.81e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.3e-07 5 4.31e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.7e-07 5 4.71e-07 0 5e-07 0 
+ 5.01e-07 5 5.3e-07 5 5.31e-07 0 5.6e-07 0 
+ 5.61e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.3e-07 5 6.31e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.9e-07 5 6.91e-07 0 7e-07 0 
+ 7.01e-07 5 7.1e-07 5 7.11e-07 0 7.3e-07 0 
+ 7.31e-07 5 7.4e-07 5 7.41e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.7e-07 5 7.71e-07 0 7.9e-07 0 
+ 7.91e-07 5 8e-07 5 8.01e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.5e-07 5 8.51e-07 0 8.8e-07 0 
+ 8.81e-07 5 9e-07 5 9.01e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.05e-06 5 )
Vaa2 565 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 7e-08 5 7.1e-08 0 8e-08 0 
+ 8.1e-08 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.4e-07 5 2.41e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.1e-07 5 3.11e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.3e-07 5 3.31e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 3.9e-07 0 
+ 3.91e-07 5 4e-07 5 4.01e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.7e-07 5 4.71e-07 0 4.8e-07 0 
+ 4.81e-07 5 4.9e-07 5 4.91e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.3e-07 5 5.31e-07 0 5.6e-07 0 
+ 5.61e-07 5 6e-07 5 6.01e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.5e-07 5 6.51e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.8e-07 5 6.81e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.8e-07 5 7.81e-07 0 7.9e-07 0 
+ 7.91e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 9.1e-07 5 9.11e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.5e-07 5 9.51e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.02e-06 5 )
Vaa3 598 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 6e-08 0 6.1e-08 5 1.1e-07 5 
+ 1.11e-07 0 1.2e-07 0 1.21e-07 5 1.3e-07 5 
+ 1.31e-07 0 1.4e-07 0 1.41e-07 5 1.8e-07 5 
+ 1.81e-07 0 2.1e-07 0 2.11e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.5e-07 0 2.51e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.5e-07 0 3.51e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.8e-07 0 3.81e-07 5 4e-07 5 
+ 4.01e-07 0 4.3e-07 0 4.31e-07 5 4.6e-07 5 
+ 4.61e-07 0 4.8e-07 0 4.81e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.1e-07 0 5.11e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.6e-07 0 5.61e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6.1e-07 0 6.11e-07 5 6.2e-07 5 
+ 6.21e-07 0 6.3e-07 0 6.31e-07 5 6.4e-07 5 
+ 6.41e-07 0 6.5e-07 0 6.51e-07 5 6.9e-07 5 
+ 6.91e-07 0 7.3e-07 0 7.31e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.8e-07 0 7.81e-07 5 8e-07 5 
+ 8.01e-07 0 8.3e-07 0 8.31e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.7e-07 0 8.71e-07 5 8.8e-07 5 
+ 8.81e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.2e-07 0 9.21e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.4e-07 0 9.41e-07 5 9.7e-07 5 
+ 9.71e-07 0 1e-06 0 1.01e-06 0 )
Vaa4 631 0 pwl (0 5 1e-08 5 1.1e-08 0 3e-08 0 
+ 3.1e-08 5 7e-08 5 7.1e-08 0 8e-08 0 
+ 8.1e-08 5 9e-08 5 9.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.4e-07 5 1.41e-07 0 1.7e-07 0 
+ 1.71e-07 5 1.9e-07 5 1.91e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.3e-07 5 2.31e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.6e-07 5 2.61e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.1e-07 5 3.11e-07 0 3.5e-07 0 
+ 3.51e-07 5 3.6e-07 5 3.61e-07 0 3.7e-07 0 
+ 3.71e-07 5 3.8e-07 5 3.81e-07 0 3.9e-07 0 
+ 3.91e-07 5 4e-07 5 4.01e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.5e-07 5 4.51e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.1e-07 5 5.11e-07 0 5.2e-07 0 
+ 5.21e-07 5 5.4e-07 5 5.41e-07 0 5.5e-07 0 
+ 5.51e-07 5 5.6e-07 5 5.61e-07 0 5.8e-07 0 
+ 5.81e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.5e-07 5 6.51e-07 0 6.7e-07 0 
+ 6.71e-07 5 7.1e-07 5 7.11e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.8e-07 5 7.81e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.5e-07 5 8.51e-07 0 8.7e-07 0 
+ 8.71e-07 5 9e-07 5 9.01e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.4e-07 5 9.41e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.6e-07 5 9.61e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 1e-06 0 
+ 1.001e-06 5 1.01e-06 5 )
Vaa5 664 0 pwl (0 5 1e-08 5 1.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 6e-08 5 6.1e-08 0 7e-08 0 
+ 7.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.4e-07 5 1.41e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.6e-07 5 1.61e-07 0 1.9e-07 0 
+ 1.91e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.2e-07 5 2.21e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.7e-07 5 2.71e-07 0 2.8e-07 0 
+ 2.81e-07 5 3.1e-07 5 3.11e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.3e-07 5 3.31e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.8e-07 0 
+ 3.81e-07 5 4.1e-07 5 4.11e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.3e-07 5 4.31e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.9e-07 5 4.91e-07 0 5e-07 0 
+ 5.01e-07 5 5.1e-07 5 5.11e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.5e-07 5 5.51e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.9e-07 5 5.91e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.4e-07 5 6.41e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.6e-07 5 7.61e-07 0 7.8e-07 0 
+ 7.81e-07 5 7.9e-07 5 7.91e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.6e-07 5 8.61e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.8e-07 5 8.81e-07 0 9e-07 0 
+ 9.01e-07 5 9.1e-07 5 9.11e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vaa6 697 0 pwl (0 5 2e-08 5 2.1e-08 0 4e-08 0 
+ 4.1e-08 5 6e-08 5 6.1e-08 0 9e-08 0 
+ 9.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.3e-07 5 1.31e-07 0 1.8e-07 0 
+ 1.81e-07 5 1.9e-07 5 1.91e-07 0 2e-07 0 
+ 2.01e-07 5 2.1e-07 5 2.11e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.6e-07 5 2.61e-07 0 3e-07 0 
+ 3.01e-07 5 3.1e-07 5 3.11e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.9e-07 0 
+ 3.91e-07 5 4e-07 5 4.01e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.3e-07 5 4.31e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.5e-07 5 4.51e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.8e-07 5 5.81e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.7e-07 5 6.71e-07 0 6.8e-07 0 
+ 6.81e-07 5 6.9e-07 5 6.91e-07 0 7e-07 0 
+ 7.01e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.3e-07 5 7.31e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.6e-07 5 7.61e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.9e-07 5 7.91e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.5e-07 5 8.51e-07 0 8.6e-07 0 
+ 8.61e-07 5 8.9e-07 5 8.91e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.4e-07 0 
+ 9.41e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 1e-06 5 )
Vaa7 730 0 pwl (0 0 3e-08 0 3.1e-08 5 4e-08 5 
+ 4.1e-08 0 7e-08 0 7.1e-08 5 8e-08 5 
+ 8.1e-08 0 1e-07 0 1.01e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.7e-07 5 
+ 1.71e-07 0 1.9e-07 0 1.91e-07 5 2e-07 5 
+ 2.01e-07 0 2.1e-07 0 2.11e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.8e-07 5 
+ 2.81e-07 0 3.4e-07 0 3.41e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.9e-07 0 3.91e-07 5 4e-07 5 
+ 4.01e-07 0 4.1e-07 0 4.11e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.4e-07 0 4.41e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.7e-07 0 4.71e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.6e-07 0 5.61e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.6e-07 0 6.61e-07 5 6.8e-07 5 
+ 6.81e-07 0 7.1e-07 0 7.11e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.8e-07 0 7.81e-07 5 8e-07 5 
+ 8.01e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.4e-07 5 
+ 8.41e-07 0 9.1e-07 0 9.11e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 1.03e-06 0 )
Vaa8 763 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 5e-08 5 5.1e-08 0 6e-08 0 
+ 6.1e-08 5 7e-08 5 7.1e-08 0 8e-08 0 
+ 8.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.5e-07 5 1.51e-07 0 1.9e-07 0 
+ 1.91e-07 5 2.1e-07 5 2.11e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.9e-07 5 2.91e-07 0 3.2e-07 0 
+ 3.21e-07 5 4.1e-07 5 4.11e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.3e-07 5 4.31e-07 0 4.4e-07 0 
+ 4.41e-07 5 5.1e-07 5 5.11e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.9e-07 5 5.91e-07 0 6e-07 0 
+ 6.01e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.5e-07 5 7.51e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.9e-07 5 7.91e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.6e-07 5 8.61e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9.1e-07 0 
+ 9.11e-07 5 9.4e-07 5 9.41e-07 0 9.6e-07 0 
+ 9.61e-07 5 1e-06 5 1.02e-06 5 )
Vaa9 796 0 pwl (0 0 3e-08 0 3.1e-08 5 5e-08 5 
+ 5.1e-08 0 6e-08 0 6.1e-08 5 7e-08 5 
+ 7.1e-08 0 9e-08 0 9.1e-08 5 1.4e-07 5 
+ 1.41e-07 0 1.6e-07 0 1.61e-07 5 1.9e-07 5 
+ 1.91e-07 0 2e-07 0 2.01e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 3.1e-07 0 3.11e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.3e-07 0 3.31e-07 5 3.4e-07 5 
+ 3.41e-07 0 3.5e-07 0 3.51e-07 5 3.8e-07 5 
+ 3.81e-07 0 4.7e-07 0 4.71e-07 5 4.8e-07 5 
+ 4.81e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.8e-07 0 5.81e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.4e-07 5 
+ 6.41e-07 0 6.5e-07 0 6.51e-07 5 6.7e-07 5 
+ 6.71e-07 0 6.8e-07 0 6.81e-07 5 7e-07 5 
+ 7.01e-07 0 7.1e-07 0 7.11e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.9e-07 5 
+ 7.91e-07 0 8e-07 0 8.01e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.6e-07 0 8.61e-07 5 8.7e-07 5 
+ 8.71e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 9.4e-07 5 
+ 9.41e-07 0 9.6e-07 0 9.61e-07 5 9.7e-07 5 
+ 9.71e-07 0 9.8e-07 0 9.81e-07 5 9.9e-07 5 
+ 9.91e-07 0 1e-06 0 )
Vaa10 829 0 pwl (0 5 4e-08 5 4.1e-08 0 6e-08 0 
+ 6.1e-08 5 7e-08 5 7.1e-08 0 8e-08 0 
+ 8.1e-08 5 9e-08 5 9.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.8e-07 0 
+ 1.81e-07 5 1.9e-07 5 1.91e-07 0 2e-07 0 
+ 2.01e-07 5 2.2e-07 5 2.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.6e-07 5 2.61e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.5e-07 0 
+ 3.51e-07 5 3.6e-07 5 3.61e-07 0 3.7e-07 0 
+ 3.71e-07 5 4e-07 5 4.01e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.3e-07 5 4.31e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.8e-07 5 4.81e-07 0 5e-07 0 
+ 5.01e-07 5 5.1e-07 5 5.11e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.7e-07 5 5.71e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.7e-07 5 6.71e-07 0 6.9e-07 0 
+ 6.91e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.5e-07 5 7.51e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.9e-07 5 7.91e-07 0 8e-07 0 
+ 8.01e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.04e-06 5 )
Vaa11 862 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 4e-08 0 4.1e-08 5 5e-08 5 
+ 5.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1e-07 0 1.01e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.7e-07 5 
+ 1.71e-07 0 1.8e-07 0 1.81e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.2e-07 0 2.21e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.6e-07 0 2.61e-07 5 2.7e-07 5 
+ 2.71e-07 0 3.2e-07 0 3.21e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.4e-07 0 3.41e-07 5 3.7e-07 5 
+ 3.71e-07 0 3.9e-07 0 3.91e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.7e-07 0 4.71e-07 5 5e-07 5 
+ 5.01e-07 0 5.1e-07 0 5.11e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.7e-07 0 5.71e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 7.2e-07 0 7.21e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.5e-07 0 7.51e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.9e-07 0 7.91e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.8e-07 0 8.81e-07 5 8.9e-07 5 
+ 8.91e-07 0 9.1e-07 0 9.11e-07 5 9.2e-07 5 
+ 9.21e-07 0 1e-06 0 1.01e-06 0 )
Vaa12 895 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 6e-08 5 
+ 6.1e-08 0 7e-08 0 7.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1.3e-07 5 
+ 1.31e-07 0 1.5e-07 0 1.51e-07 5 1.7e-07 5 
+ 1.71e-07 0 2e-07 0 2.01e-07 5 2.1e-07 5 
+ 2.11e-07 0 2.2e-07 0 2.21e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.9e-07 0 2.91e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.3e-07 0 3.31e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.8e-07 0 3.81e-07 5 4e-07 5 
+ 4.01e-07 0 4.2e-07 0 4.21e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.5e-07 0 5.51e-07 5 5.7e-07 5 
+ 5.71e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.3e-07 0 6.31e-07 5 6.4e-07 5 
+ 6.41e-07 0 6.5e-07 0 6.51e-07 5 7.1e-07 5 
+ 7.11e-07 0 7.2e-07 0 7.21e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.6e-07 0 8.61e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 8.9e-07 5 
+ 8.91e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 9.4e-07 5 
+ 9.41e-07 0 9.5e-07 0 9.51e-07 5 9.6e-07 5 
+ 9.61e-07 0 1e-06 0 1.01e-06 0 )
Vaa13 928 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 4e-08 0 4.1e-08 5 5e-08 5 
+ 5.1e-08 0 6e-08 0 6.1e-08 5 9e-08 5 
+ 9.1e-08 0 1e-07 0 1.01e-07 5 1.1e-07 5 
+ 1.11e-07 0 1.2e-07 0 1.21e-07 5 1.3e-07 5 
+ 1.31e-07 0 1.8e-07 0 1.81e-07 5 1.9e-07 5 
+ 1.91e-07 0 2e-07 0 2.01e-07 5 2.1e-07 5 
+ 2.11e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.7e-07 0 2.71e-07 5 2.8e-07 5 
+ 2.81e-07 0 3e-07 0 3.01e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.3e-07 0 3.31e-07 5 3.4e-07 5 
+ 3.41e-07 0 3.6e-07 0 3.61e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.5e-07 0 4.51e-07 5 4.6e-07 5 
+ 4.61e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.6e-07 0 5.61e-07 5 6e-07 5 
+ 6.01e-07 0 6.3e-07 0 6.31e-07 5 6.7e-07 5 
+ 6.71e-07 0 6.8e-07 0 6.81e-07 5 6.9e-07 5 
+ 6.91e-07 0 7.1e-07 0 7.11e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.4e-07 0 8.41e-07 5 8.6e-07 5 
+ 8.61e-07 0 8.9e-07 0 8.91e-07 5 9e-07 5 
+ 9.01e-07 0 9.2e-07 0 9.21e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.7e-07 0 9.71e-07 5 1e-06 5 
+ 1.001e-06 0 1.01e-06 0 )
Vaa14 961 0 pwl (0 0 1e-08 0 1.1e-08 5 6e-08 5 
+ 6.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.2e-07 0 1.21e-07 5 1.3e-07 5 
+ 1.31e-07 0 1.5e-07 0 1.51e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.9e-07 0 1.91e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.5e-07 0 2.51e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.8e-07 0 2.81e-07 5 3e-07 5 
+ 3.01e-07 0 3.1e-07 0 3.11e-07 5 3.7e-07 5 
+ 3.71e-07 0 3.8e-07 0 3.81e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.5e-07 0 5.51e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6e-07 0 6.01e-07 5 6.2e-07 5 
+ 6.21e-07 0 6.4e-07 0 6.41e-07 5 6.5e-07 5 
+ 6.51e-07 0 6.6e-07 0 6.61e-07 5 6.8e-07 5 
+ 6.81e-07 0 6.9e-07 0 6.91e-07 5 7e-07 5 
+ 7.01e-07 0 7.1e-07 0 7.11e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.5e-07 0 7.51e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.6e-07 0 8.61e-07 5 8.7e-07 5 
+ 8.71e-07 0 9e-07 0 9.01e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.3e-07 0 9.31e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 1.01e-06 0 )
Vaa15 994 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 3e-08 0 3.1e-08 5 4e-08 5 
+ 4.1e-08 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.5e-07 5 
+ 1.51e-07 0 1.7e-07 0 1.71e-07 5 1.9e-07 5 
+ 1.91e-07 0 2e-07 0 2.01e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.4e-07 0 2.41e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.6e-07 0 2.61e-07 5 2.7e-07 5 
+ 2.71e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.1e-07 0 3.11e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.4e-07 0 3.41e-07 5 3.5e-07 5 
+ 3.51e-07 0 4e-07 0 4.01e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.4e-07 0 4.41e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 4.9e-07 5 
+ 4.91e-07 0 5e-07 0 5.01e-07 5 5.1e-07 5 
+ 5.11e-07 0 5.2e-07 0 5.21e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.5e-07 0 5.51e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.8e-07 0 5.81e-07 5 6e-07 5 
+ 6.01e-07 0 6.1e-07 0 6.11e-07 5 6.2e-07 5 
+ 6.21e-07 0 6.4e-07 0 6.41e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.7e-07 0 6.71e-07 5 7.1e-07 5 
+ 7.11e-07 0 7.2e-07 0 7.21e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8e-07 5 
+ 8.01e-07 0 8.1e-07 0 8.11e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.8e-07 0 8.81e-07 5 8.9e-07 5 
+ 8.91e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.8e-07 0 9.81e-07 5 1e-06 5 
+ 1.001e-06 0 )
Vaa16 1027 0 pwl (0 5 3e-08 5 3.1e-08 0 7e-08 0 
+ 7.1e-08 5 8e-08 5 8.1e-08 0 1.5e-07 0 
+ 1.51e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.4e-07 5 2.41e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.7e-07 5 2.71e-07 0 2.8e-07 0 
+ 2.81e-07 5 3e-07 5 3.01e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.2e-07 5 3.21e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.8e-07 0 
+ 3.81e-07 5 4e-07 5 4.01e-07 0 4.2e-07 0 
+ 4.21e-07 5 4.4e-07 5 4.41e-07 0 4.6e-07 0 
+ 4.61e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.8e-07 5 5.81e-07 0 6e-07 0 
+ 6.01e-07 5 6.1e-07 5 6.11e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.8e-07 5 6.81e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.3e-07 5 7.31e-07 0 7.8e-07 0 
+ 7.81e-07 5 8.1e-07 5 8.11e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.4e-07 5 8.41e-07 0 8.5e-07 0 
+ 8.51e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9e-07 0 
+ 9.01e-07 5 9.2e-07 5 9.21e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.6e-07 5 9.61e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.03e-06 5 )
Vbb1 533 0 pwl (0 5 3e-08 5 3.1e-08 0 4e-08 0 
+ 4.1e-08 5 5e-08 5 5.1e-08 0 9e-08 0 
+ 9.1e-08 5 1e-07 5 1.01e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 2.4e-07 5 2.41e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.8e-07 5 2.81e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.2e-07 5 3.21e-07 0 3.3e-07 0 
+ 3.31e-07 5 3.4e-07 5 3.41e-07 0 3.7e-07 0 
+ 3.71e-07 5 3.8e-07 5 3.81e-07 0 4e-07 0 
+ 4.01e-07 5 4.2e-07 5 4.21e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.4e-07 5 4.41e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.6e-07 5 4.61e-07 0 4.7e-07 0 
+ 4.71e-07 5 4.8e-07 5 4.81e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.4e-07 5 5.41e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.9e-07 5 5.91e-07 0 6e-07 0 
+ 6.01e-07 5 6.1e-07 5 6.11e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.4e-07 5 6.41e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.9e-07 5 6.91e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.9e-07 5 7.91e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.7e-07 5 8.71e-07 0 9e-07 0 
+ 9.01e-07 5 9.1e-07 5 9.11e-07 0 9.9e-07 0 
+ 9.91e-07 5 1e-06 5 1.03e-06 5 )
Vbb2 566 0 pwl (0 5 3e-08 5 3.1e-08 0 6e-08 0 
+ 6.1e-08 5 8e-08 5 8.1e-08 0 9e-08 0 
+ 9.1e-08 5 1e-07 5 1.01e-07 0 1.1e-07 0 
+ 1.11e-07 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.5e-07 5 1.51e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.7e-07 5 1.71e-07 0 1.8e-07 0 
+ 1.81e-07 5 2.2e-07 5 2.21e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.3e-07 5 3.31e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.7e-07 5 3.71e-07 0 4e-07 0 
+ 4.01e-07 5 4.2e-07 5 4.21e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.6e-07 5 4.61e-07 0 4.7e-07 0 
+ 4.71e-07 5 4.8e-07 5 4.81e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.3e-07 5 5.31e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.9e-07 5 5.91e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.3e-07 5 6.31e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.8e-07 5 6.81e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.3e-07 5 7.31e-07 0 7.6e-07 0 
+ 7.61e-07 5 7.7e-07 5 7.71e-07 0 7.9e-07 0 
+ 7.91e-07 5 8e-07 5 8.01e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.4e-07 5 8.41e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.6e-07 5 9.61e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vbb3 599 0 pwl (0 0 2e-08 0 2.1e-08 5 3e-08 5 
+ 3.1e-08 0 6e-08 0 6.1e-08 5 7e-08 5 
+ 7.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.5e-07 5 
+ 1.51e-07 0 1.6e-07 0 1.61e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.3e-07 0 2.31e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.6e-07 0 2.61e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.4e-07 0 3.41e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 3.9e-07 5 
+ 3.91e-07 0 4e-07 0 4.01e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.3e-07 0 4.31e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 4.7e-07 5 
+ 4.71e-07 0 5e-07 0 5.01e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.4e-07 0 5.41e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.6e-07 0 5.61e-07 5 5.8e-07 5 
+ 5.81e-07 0 5.9e-07 0 5.91e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.4e-07 0 6.41e-07 5 6.5e-07 5 
+ 6.51e-07 0 6.6e-07 0 6.61e-07 5 6.7e-07 5 
+ 6.71e-07 0 6.9e-07 0 6.91e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.4e-07 0 7.41e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.3e-07 5 
+ 8.31e-07 0 8.9e-07 0 8.91e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 1e-06 5 
+ 1.001e-06 0 1.02e-06 0 )
Vbb4 632 0 pwl (0 5 1e-08 5 1.1e-08 0 2e-08 0 
+ 2.1e-08 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 6e-08 5 6.1e-08 0 7e-08 0 
+ 7.1e-08 5 8e-08 5 8.1e-08 0 1.1e-07 0 
+ 1.11e-07 5 1.3e-07 5 1.31e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.9e-07 5 1.91e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.2e-07 5 2.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3e-07 5 3.01e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.3e-07 5 3.31e-07 0 3.8e-07 0 
+ 3.81e-07 5 3.9e-07 5 3.91e-07 0 4e-07 0 
+ 4.01e-07 5 4.4e-07 5 4.41e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.7e-07 5 4.71e-07 0 4.9e-07 0 
+ 4.91e-07 5 5e-07 5 5.01e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 6.3e-07 5 6.31e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 6.7e-07 0 
+ 6.71e-07 5 6.9e-07 5 6.91e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.3e-07 5 7.31e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.8e-07 5 7.81e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.5e-07 0 
+ 8.51e-07 5 8.7e-07 5 8.71e-07 0 8.8e-07 0 
+ 8.81e-07 5 8.9e-07 5 8.91e-07 0 9e-07 0 
+ 9.01e-07 5 9.6e-07 5 9.61e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vbb5 665 0 pwl (0 0 2e-08 0 2.1e-08 5 4e-08 5 
+ 4.1e-08 0 6e-08 0 6.1e-08 5 7e-08 5 
+ 7.1e-08 0 8e-08 0 8.1e-08 5 9e-08 5 
+ 9.1e-08 0 1.1e-07 0 1.11e-07 5 1.5e-07 5 
+ 1.51e-07 0 1.6e-07 0 1.61e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.4e-07 0 2.41e-07 5 2.5e-07 5 
+ 2.51e-07 0 2.7e-07 0 2.71e-07 5 2.9e-07 5 
+ 2.91e-07 0 3.1e-07 0 3.11e-07 5 3.3e-07 5 
+ 3.31e-07 0 3.5e-07 0 3.51e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 4.2e-07 5 
+ 4.21e-07 0 4.3e-07 0 4.31e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.7e-07 0 4.71e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.1e-07 0 5.11e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6.3e-07 0 6.31e-07 5 6.4e-07 5 
+ 6.41e-07 0 6.5e-07 0 6.51e-07 5 6.7e-07 5 
+ 6.71e-07 0 6.8e-07 0 6.81e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.6e-07 0 7.61e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.8e-07 0 7.81e-07 5 8e-07 5 
+ 8.01e-07 0 8.1e-07 0 8.11e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.4e-07 0 8.41e-07 5 8.6e-07 5 
+ 8.61e-07 0 8.9e-07 0 8.91e-07 5 9e-07 5 
+ 9.01e-07 0 9.2e-07 0 9.21e-07 5 9.3e-07 5 
+ 9.31e-07 0 9.4e-07 0 9.41e-07 5 9.7e-07 5 
+ 9.71e-07 0 1e-06 0 )
Vbb6 698 0 pwl (0 5 4e-08 5 4.1e-08 0 5e-08 0 
+ 5.1e-08 5 7e-08 5 7.1e-08 0 9e-08 0 
+ 9.1e-08 5 1.3e-07 5 1.31e-07 0 1.4e-07 0 
+ 1.41e-07 5 1.6e-07 5 1.61e-07 0 1.7e-07 0 
+ 1.71e-07 5 2e-07 5 2.01e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.5e-07 5 2.51e-07 0 2.6e-07 0 
+ 2.61e-07 5 2.8e-07 5 2.81e-07 0 3e-07 0 
+ 3.01e-07 5 3.6e-07 5 3.61e-07 0 3.8e-07 0 
+ 3.81e-07 5 3.9e-07 5 3.91e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.2e-07 5 4.21e-07 0 4.4e-07 0 
+ 4.41e-07 5 4.6e-07 5 4.61e-07 0 5e-07 0 
+ 5.01e-07 5 5.2e-07 5 5.21e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.7e-07 5 5.71e-07 0 5.8e-07 0 
+ 5.81e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.9e-07 5 6.91e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.3e-07 5 7.31e-07 0 7.4e-07 0 
+ 7.41e-07 5 7.5e-07 5 7.51e-07 0 7.9e-07 0 
+ 7.91e-07 5 8.3e-07 5 8.31e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.6e-07 5 8.61e-07 0 8.9e-07 0 
+ 8.91e-07 5 9e-07 5 9.01e-07 0 9.3e-07 0 
+ 9.31e-07 5 9.5e-07 5 9.51e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vbb7 731 0 pwl (0 5 1e-08 5 1.1e-08 0 4e-08 0 
+ 4.1e-08 5 5e-08 5 5.1e-08 0 6e-08 0 
+ 6.1e-08 5 7e-08 5 7.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.3e-07 0 
+ 1.31e-07 5 1.5e-07 5 1.51e-07 0 1.8e-07 0 
+ 1.81e-07 5 2e-07 5 2.01e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.2e-07 5 2.21e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.7e-07 5 2.71e-07 0 2.8e-07 0 
+ 2.81e-07 5 2.9e-07 5 2.91e-07 0 3.1e-07 0 
+ 3.11e-07 5 3.7e-07 5 3.71e-07 0 4e-07 0 
+ 4.01e-07 5 4.3e-07 5 4.31e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.9e-07 5 4.91e-07 0 5.1e-07 0 
+ 5.11e-07 5 5.3e-07 5 5.31e-07 0 5.5e-07 0 
+ 5.51e-07 5 5.6e-07 5 5.61e-07 0 5.8e-07 0 
+ 5.81e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 7e-07 5 7.01e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.6e-07 5 7.61e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.8e-07 5 7.81e-07 0 8e-07 0 
+ 8.01e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 9.3e-07 5 9.31e-07 0 9.7e-07 0 
+ 9.71e-07 5 1e-06 5 )
Vbb8 764 0 pwl (0 5 3e-08 5 3.1e-08 0 4e-08 0 
+ 4.1e-08 5 5e-08 5 5.1e-08 0 7e-08 0 
+ 7.1e-08 5 8e-08 5 8.1e-08 0 9e-08 0 
+ 9.1e-08 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.3e-07 5 1.31e-07 0 1.5e-07 0 
+ 1.51e-07 5 1.8e-07 5 1.81e-07 0 2e-07 0 
+ 2.01e-07 5 2.5e-07 5 2.51e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.3e-07 5 3.31e-07 0 3.9e-07 0 
+ 3.91e-07 5 4.1e-07 5 4.11e-07 0 4.5e-07 0 
+ 4.51e-07 5 4.7e-07 5 4.71e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.1e-07 5 5.11e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.5e-07 5 5.51e-07 0 5.6e-07 0 
+ 5.61e-07 5 5.7e-07 5 5.71e-07 0 5.8e-07 0 
+ 5.81e-07 5 6e-07 5 6.01e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.2e-07 5 6.21e-07 0 6.3e-07 0 
+ 6.31e-07 5 6.4e-07 5 6.41e-07 0 6.5e-07 0 
+ 6.51e-07 5 6.6e-07 5 6.61e-07 0 6.7e-07 0 
+ 6.71e-07 5 7e-07 5 7.01e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.3e-07 5 7.31e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.9e-07 5 7.91e-07 0 8.1e-07 0 
+ 8.11e-07 5 8.2e-07 5 8.21e-07 0 8.3e-07 0 
+ 8.31e-07 5 8.4e-07 5 8.41e-07 0 8.7e-07 0 
+ 8.71e-07 5 8.8e-07 5 8.81e-07 0 9.2e-07 0 
+ 9.21e-07 5 9.3e-07 5 9.31e-07 0 9.5e-07 0 
+ 9.51e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 1.03e-06 5 )
Vbb9 797 0 pwl (0 0 2e-08 0 2.1e-08 5 4e-08 5 
+ 4.1e-08 0 5e-08 0 5.1e-08 5 6e-08 5 
+ 6.1e-08 0 7e-08 0 7.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.8e-07 0 1.81e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.2e-07 0 2.21e-07 5 2.4e-07 5 
+ 2.41e-07 0 2.6e-07 0 2.61e-07 5 2.8e-07 5 
+ 2.81e-07 0 3e-07 0 3.01e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.4e-07 0 3.41e-07 5 3.7e-07 5 
+ 3.71e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4.2e-07 0 4.21e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.8e-07 0 4.81e-07 5 5e-07 5 
+ 5.01e-07 0 5.1e-07 0 5.11e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.6e-07 0 5.61e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 6e-07 5 
+ 6.01e-07 0 6.1e-07 0 6.11e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.4e-07 0 6.41e-07 5 6.5e-07 5 
+ 6.51e-07 0 6.7e-07 0 6.71e-07 5 6.8e-07 5 
+ 6.81e-07 0 7e-07 0 7.01e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.5e-07 0 7.51e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.8e-07 5 
+ 7.81e-07 0 7.9e-07 0 7.91e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.6e-07 0 8.61e-07 5 8.8e-07 5 
+ 8.81e-07 0 8.9e-07 0 8.91e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 9.4e-07 5 
+ 9.41e-07 0 1e-06 0 )
Vbb10 830 0 pwl (0 0 2e-08 0 2.1e-08 5 8e-08 5 
+ 8.1e-08 0 1.2e-07 0 1.21e-07 5 1.7e-07 5 
+ 1.71e-07 0 1.8e-07 0 1.81e-07 5 1.9e-07 5 
+ 1.91e-07 0 2e-07 0 2.01e-07 5 2.1e-07 5 
+ 2.11e-07 0 2.2e-07 0 2.21e-07 5 2.3e-07 5 
+ 2.31e-07 0 2.8e-07 0 2.81e-07 5 2.9e-07 5 
+ 2.91e-07 0 3e-07 0 3.01e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.3e-07 0 3.31e-07 5 3.4e-07 5 
+ 3.41e-07 0 3.5e-07 0 3.51e-07 5 3.8e-07 5 
+ 3.81e-07 0 4.6e-07 0 4.61e-07 5 5e-07 5 
+ 5.01e-07 0 5.4e-07 0 5.41e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 5.9e-07 5 
+ 5.91e-07 0 6e-07 0 6.01e-07 5 6.1e-07 5 
+ 6.11e-07 0 6.4e-07 0 6.41e-07 5 6.5e-07 5 
+ 6.51e-07 0 6.7e-07 0 6.71e-07 5 6.9e-07 5 
+ 6.91e-07 0 7.2e-07 0 7.21e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.4e-07 0 7.41e-07 5 7.6e-07 5 
+ 7.61e-07 0 7.7e-07 0 7.71e-07 5 7.9e-07 5 
+ 7.91e-07 0 8e-07 0 8.01e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.3e-07 0 8.31e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.5e-07 0 8.51e-07 5 9e-07 5 
+ 9.01e-07 0 9.1e-07 0 9.11e-07 5 9.2e-07 5 
+ 9.21e-07 0 9.3e-07 0 9.31e-07 5 9.4e-07 5 
+ 9.41e-07 0 9.5e-07 0 9.51e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 1.02e-06 0 )
Vbb11 863 0 pwl (0 0 1e-08 0 1.1e-08 5 6e-08 5 
+ 6.1e-08 0 7e-08 0 7.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 1.7e-07 0 1.71e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.3e-07 0 2.31e-07 5 2.8e-07 5 
+ 2.81e-07 0 2.9e-07 0 2.91e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.8e-07 0 3.81e-07 5 4e-07 5 
+ 4.01e-07 0 4.2e-07 0 4.21e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.7e-07 0 4.71e-07 5 4.8e-07 5 
+ 4.81e-07 0 4.9e-07 0 4.91e-07 5 5e-07 5 
+ 5.01e-07 0 5.2e-07 0 5.21e-07 5 5.3e-07 5 
+ 5.31e-07 0 5.4e-07 0 5.41e-07 5 5.6e-07 5 
+ 5.61e-07 0 5.7e-07 0 5.71e-07 5 5.8e-07 5 
+ 5.81e-07 0 5.9e-07 0 5.91e-07 5 6e-07 5 
+ 6.01e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.5e-07 0 6.51e-07 5 6.8e-07 5 
+ 6.81e-07 0 6.9e-07 0 6.91e-07 5 7.1e-07 5 
+ 7.11e-07 0 7.4e-07 0 7.41e-07 5 7.7e-07 5 
+ 7.71e-07 0 7.8e-07 0 7.81e-07 5 8.5e-07 5 
+ 8.51e-07 0 8.6e-07 0 8.61e-07 5 8.8e-07 5 
+ 8.81e-07 0 9e-07 0 9.01e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.5e-07 0 9.51e-07 5 9.6e-07 5 
+ 9.61e-07 0 9.7e-07 0 9.71e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 )
Vbb12 896 0 pwl (0 5 2e-08 5 2.1e-08 0 3e-08 0 
+ 3.1e-08 5 4e-08 5 4.1e-08 0 6e-08 0 
+ 6.1e-08 5 8e-08 5 8.1e-08 0 9e-08 0 
+ 9.1e-08 5 1.4e-07 5 1.41e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.8e-07 5 1.81e-07 0 2.1e-07 0 
+ 2.11e-07 5 2.2e-07 5 2.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 2.6e-07 5 2.61e-07 0 2.7e-07 0 
+ 2.71e-07 5 2.8e-07 5 2.81e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.4e-07 5 3.41e-07 0 3.6e-07 0 
+ 3.61e-07 5 3.8e-07 5 3.81e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.2e-07 5 4.21e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.6e-07 5 4.61e-07 0 4.8e-07 0 
+ 4.81e-07 5 4.9e-07 5 4.91e-07 0 5e-07 0 
+ 5.01e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.6e-07 5 5.61e-07 0 5.7e-07 0 
+ 5.71e-07 5 6.1e-07 5 6.11e-07 0 6.2e-07 0 
+ 6.21e-07 5 6.3e-07 5 6.31e-07 0 6.4e-07 0 
+ 6.41e-07 5 6.8e-07 5 6.81e-07 0 6.9e-07 0 
+ 6.91e-07 5 7.1e-07 5 7.11e-07 0 7.3e-07 0 
+ 7.31e-07 5 7.4e-07 5 7.41e-07 0 7.7e-07 0 
+ 7.71e-07 5 7.9e-07 5 7.91e-07 0 8e-07 0 
+ 8.01e-07 5 8.1e-07 5 8.11e-07 0 8.2e-07 0 
+ 8.21e-07 5 8.3e-07 5 8.31e-07 0 8.6e-07 0 
+ 8.61e-07 5 8.7e-07 5 8.71e-07 0 8.9e-07 0 
+ 8.91e-07 5 9.3e-07 5 9.31e-07 0 9.6e-07 0 
+ 9.61e-07 5 1e-06 5 )
Vbb13 929 0 pwl (0 0 1e-08 0 1.1e-08 5 2e-08 5 
+ 2.1e-08 0 4e-08 0 4.1e-08 5 5e-08 5 
+ 5.1e-08 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 9e-08 0 9.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.2e-07 0 1.21e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.5e-07 0 1.51e-07 5 1.6e-07 5 
+ 1.61e-07 0 2e-07 0 2.01e-07 5 2.2e-07 5 
+ 2.21e-07 0 2.7e-07 0 2.71e-07 5 2.8e-07 5 
+ 2.81e-07 0 3e-07 0 3.01e-07 5 3.1e-07 5 
+ 3.11e-07 0 3.2e-07 0 3.21e-07 5 3.5e-07 5 
+ 3.51e-07 0 3.8e-07 0 3.81e-07 5 3.9e-07 5 
+ 3.91e-07 0 4.4e-07 0 4.41e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 5e-07 5 
+ 5.01e-07 0 5.1e-07 0 5.11e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.4e-07 0 5.41e-07 5 5.5e-07 5 
+ 5.51e-07 0 5.6e-07 0 5.61e-07 5 5.7e-07 5 
+ 5.71e-07 0 5.8e-07 0 5.81e-07 5 6.2e-07 5 
+ 6.21e-07 0 6.8e-07 0 6.81e-07 5 6.9e-07 5 
+ 6.91e-07 0 7e-07 0 7.01e-07 5 7.4e-07 5 
+ 7.41e-07 0 7.6e-07 0 7.61e-07 5 7.8e-07 5 
+ 7.81e-07 0 8e-07 0 8.01e-07 5 8.1e-07 5 
+ 8.11e-07 0 8.2e-07 0 8.21e-07 5 8.4e-07 5 
+ 8.41e-07 0 8.7e-07 0 8.71e-07 5 8.8e-07 5 
+ 8.81e-07 0 9.4e-07 0 9.41e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.6e-07 0 9.61e-07 5 9.8e-07 5 
+ 9.81e-07 0 9.9e-07 0 9.91e-07 5 1e-06 5 
+ 1.001e-06 0 )
Vbb14 962 0 pwl (0 5 3e-08 5 3.1e-08 0 6e-08 0 
+ 6.1e-08 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.6e-07 5 1.61e-07 0 1.9e-07 0 
+ 1.91e-07 5 2.1e-07 5 2.11e-07 0 2.2e-07 0 
+ 2.21e-07 5 2.3e-07 5 2.31e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.6e-07 5 2.61e-07 0 2.9e-07 0 
+ 2.91e-07 5 3.1e-07 5 3.11e-07 0 3.2e-07 0 
+ 3.21e-07 5 3.5e-07 5 3.51e-07 0 3.6e-07 0 
+ 3.61e-07 5 4.1e-07 5 4.11e-07 0 4.3e-07 0 
+ 4.31e-07 5 4.6e-07 5 4.61e-07 0 4.7e-07 0 
+ 4.71e-07 5 5.2e-07 5 5.21e-07 0 5.3e-07 0 
+ 5.31e-07 5 5.4e-07 5 5.41e-07 0 5.7e-07 0 
+ 5.71e-07 5 5.9e-07 5 5.91e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.3e-07 5 6.31e-07 0 6.9e-07 0 
+ 6.91e-07 5 7e-07 5 7.01e-07 0 7.1e-07 0 
+ 7.11e-07 5 7.7e-07 5 7.71e-07 0 7.8e-07 0 
+ 7.81e-07 5 8.3e-07 5 8.31e-07 0 8.5e-07 0 
+ 8.51e-07 5 8.6e-07 5 8.61e-07 0 8.9e-07 0 
+ 8.91e-07 5 9.2e-07 5 9.21e-07 0 9.6e-07 0 
+ 9.61e-07 5 9.7e-07 5 9.71e-07 0 9.8e-07 0 
+ 9.81e-07 5 9.9e-07 5 9.91e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vbb15 995 0 pwl (0 5 1e-08 5 1.1e-08 0 3e-08 0 
+ 3.1e-08 5 5e-08 5 5.1e-08 0 7e-08 0 
+ 7.1e-08 5 8e-08 5 8.1e-08 0 1e-07 0 
+ 1.01e-07 5 1.1e-07 5 1.11e-07 0 1.2e-07 0 
+ 1.21e-07 5 1.4e-07 5 1.41e-07 0 1.6e-07 0 
+ 1.61e-07 5 1.9e-07 5 1.91e-07 0 2.3e-07 0 
+ 2.31e-07 5 2.4e-07 5 2.41e-07 0 2.5e-07 0 
+ 2.51e-07 5 2.6e-07 5 2.61e-07 0 2.7e-07 0 
+ 2.71e-07 5 2.8e-07 5 2.81e-07 0 3e-07 0 
+ 3.01e-07 5 3.1e-07 5 3.11e-07 0 3.4e-07 0 
+ 3.41e-07 5 3.5e-07 5 3.51e-07 0 4.1e-07 0 
+ 4.11e-07 5 4.5e-07 5 4.51e-07 0 4.6e-07 0 
+ 4.61e-07 5 4.7e-07 5 4.71e-07 0 4.9e-07 0 
+ 4.91e-07 5 5.1e-07 5 5.11e-07 0 5.4e-07 0 
+ 5.41e-07 5 5.7e-07 5 5.71e-07 0 5.8e-07 0 
+ 5.81e-07 5 5.9e-07 5 5.91e-07 0 6.1e-07 0 
+ 6.11e-07 5 6.2e-07 5 6.21e-07 0 6.6e-07 0 
+ 6.61e-07 5 6.7e-07 5 6.71e-07 0 6.8e-07 0 
+ 6.81e-07 5 7.1e-07 5 7.11e-07 0 7.2e-07 0 
+ 7.21e-07 5 7.4e-07 5 7.41e-07 0 7.5e-07 0 
+ 7.51e-07 5 7.6e-07 5 7.61e-07 0 7.8e-07 0 
+ 7.81e-07 5 8.1e-07 5 8.11e-07 0 8.4e-07 0 
+ 8.41e-07 5 8.7e-07 5 8.71e-07 0 8.9e-07 0 
+ 8.91e-07 5 9e-07 5 9.01e-07 0 9.7e-07 0 
+ 9.71e-07 5 9.8e-07 5 9.81e-07 0 1e-06 0 
+ 1.001e-06 5 )
Vbb16 1028 0 pwl (0 0 2e-08 0 2.1e-08 5 4e-08 5 
+ 4.1e-08 0 6e-08 0 6.1e-08 5 1e-07 5 
+ 1.01e-07 0 1.1e-07 0 1.11e-07 5 1.2e-07 5 
+ 1.21e-07 0 1.3e-07 0 1.31e-07 5 1.4e-07 5 
+ 1.41e-07 0 1.6e-07 0 1.61e-07 5 1.9e-07 5 
+ 1.91e-07 0 2.3e-07 0 2.31e-07 5 2.6e-07 5 
+ 2.61e-07 0 2.7e-07 0 2.71e-07 5 2.9e-07 5 
+ 2.91e-07 0 3e-07 0 3.01e-07 5 3.6e-07 5 
+ 3.61e-07 0 3.7e-07 0 3.71e-07 5 3.8e-07 5 
+ 3.81e-07 0 3.9e-07 0 3.91e-07 5 4.1e-07 5 
+ 4.11e-07 0 4.2e-07 0 4.21e-07 5 4.3e-07 5 
+ 4.31e-07 0 4.4e-07 0 4.41e-07 5 4.5e-07 5 
+ 4.51e-07 0 4.6e-07 0 4.61e-07 5 4.7e-07 5 
+ 4.71e-07 0 4.8e-07 0 4.81e-07 5 4.9e-07 5 
+ 4.91e-07 0 5.1e-07 0 5.11e-07 5 5.2e-07 5 
+ 5.21e-07 0 5.3e-07 0 5.31e-07 5 5.4e-07 5 
+ 5.41e-07 0 5.5e-07 0 5.51e-07 5 5.9e-07 5 
+ 5.91e-07 0 6.2e-07 0 6.21e-07 5 6.3e-07 5 
+ 6.31e-07 0 6.5e-07 0 6.51e-07 5 6.6e-07 5 
+ 6.61e-07 0 6.9e-07 0 6.91e-07 5 7e-07 5 
+ 7.01e-07 0 7.2e-07 0 7.21e-07 5 7.3e-07 5 
+ 7.31e-07 0 7.4e-07 0 7.41e-07 5 7.5e-07 5 
+ 7.51e-07 0 7.6e-07 0 7.61e-07 5 7.9e-07 5 
+ 7.91e-07 0 8e-07 0 8.01e-07 5 8.2e-07 5 
+ 8.21e-07 0 8.5e-07 0 8.51e-07 5 8.7e-07 5 
+ 8.71e-07 0 8.8e-07 0 8.81e-07 5 9.1e-07 5 
+ 9.11e-07 0 9.3e-07 0 9.31e-07 5 9.5e-07 5 
+ 9.51e-07 0 9.6e-07 0 9.61e-07 5 9.9e-07 5 
+ 9.91e-07 0 1e-06 0 )
VCIN 5 0 0 
VVDD 1 0 5
.op
*.print TRAN v(3) v(4) v(5) v(6) v(7) v(37) 
+v(38) v(7) v(39) v(40) v(70) v(71) 
+v(40) v(72) v(73) v(103) v(104) v(73) 
+v(105) v(106) v(136) v(137) v(106) v(138) 
+v(139) v(169) v(170) v(139) v(171) v(172) 
+v(202) v(203) v(172) v(204) v(205) v(235) 
+v(236) v(205) v(237) v(238) 
.options limpts=50000 itl5=50000
*.TRAN 1e-09 1e-06
.end
