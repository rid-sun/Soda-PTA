* RCA3040 - WIDEBAND AMP.
RS1 30 1 1K
RS2 31 0 1K
R1 5 3 4.8K
R2 6 3 4.8K
R3 9 3 811
R4 8 3 2.17K
R5 8 0 820
R6 2 14 1.32K
R7 2 12 4.5K
R8 2 15 1.32K
R9 16 0 5.25K
R10 17 0 5.25K
Q1 2 30 5 0 QNL
Q2 2 31 6 0 QNL
Q3 10 5 7 0 QNL
Q4 11 6 7 0 QNL
Q5 14 12 10 0 QNL
Q6 15 12 11 0 QNL
Q7 12 12 13 0 QNL
Q8 13 13 0 0 QNL
Q9 7 8 9 0 QNL
Q10 2 15 16 0 QNL
Q11 2 14 17 0 QNL
.MODEL QNL NPN BF=80 RB=100 TF=0.3NS TR=6NS CJE=3PF CJC=2PF VA=50
*.MODEL QNL NPN  BF=50 BR=1 IS=1e-14 RB=70 RC=40 VAF=50 TF=1E-10 TR=1E-8
*+              CJE=9e-13 CJC=1.5e-12 

*
VIN 1 0 SIN(0 0.1 50MEG 0.5NS 0.0)
VCC 2 0 DC 15.0
VEE 3 0 DC -15.0
*.PRINT DC V(1) V(2) V(3) V(4) V(5) V(6) V(7) V(8) V(9) V(10) V(11)
*+ V(12) V(13) V(14) V(15) V(16) V(17)
*.PRINT TRAN V(1) V(16) V(17)
*.TRAN 0.5NS 250NS
.OPTIONS LIMPTS=501
.op
.END
