* "Wide" nfet model (use nnfet for widths less than about 4u)
.model nfet nmos
+     Level=3          Uo=515          Vto=0.88      Tox=265e-10     
+     NSub=2.8e+16     Gamma=0.45      Phi=0.56
+     Ld=0.205u      Xj=0.25u     VMax=1.43e+5     Delta=0.2
+     Js=1000u     Pb=0.8          Cgso=245p      Cgdo=245p     
+     Cgbo=430p     Cj=250u      Cjsw=290p     Mjsw=0.3     
+     Fc=0           Tpg=1.0     
+     Theta=0.045     Eta=0.02     Kappa=0.3
*+     Wd=0.76u
*+     Rsh=70
     
* "Narrow" nfet model; use for widths less than about 4u:
.model nnfet nmos
+     Level=3          Uo=515          Vto=0.90      Tox=265e-10     
+     NSub=2.8e+16     Gamma=0.52      Phi=0.56
+     Ld=0.205u      Xj=0.25u     VMax=1.43e+5     Delta=0.2
+     Js=1000u     Pb=0.8          Cgso=245p      Cgdo=245p     
+     Cgbo=430p     Cj=250u      Cjsw=290p     Mjsw=0.3     
+     Fc=0           Tpg=1.0     
+     Theta=0.045     Eta=0.02     Kappa=0.3
*+     Wd=0.76u
*+     Rsh=70

* "Wide" pfet model (use npfet for widths less than 4u):
.model pfet pmos
+     Level=3          Uo=193          Vto=-0.80      Tox=265e-10     
+     NSub=2.8e+16     Gamma=0.50      Phi=0.60
+     Ld=-0.025u      Xj=0.20u     VMax=2.3e+5     Delta=0
+     Js=1000u     Pb=0.9          Cgso=245p      Cgdo=245p     
+     Cgbo=430p     Cj=720u      Cjsw=255p     Mjsw=0.3     
+      Fc=0           Tpg=-1.0
+     Theta=0.12     Eta=0.02     Kappa=10.0
*+     Wd=0.78u
*+     Rsh=150

* "Narrow" pfet model; use for widths less than 4u:
.model npfet pmos
+     Level=3          Uo=193          Vto=-1.05      Tox=265e-10     
+     NSub=2.8e+16     Gamma=0.70      Phi=0.60
+     Ld=-0.025u      Xj=0.20u     VMax=2.3e+5     Delta=0
+     Js=1000u     Pb=0.9          Cgso=245p      Cgdo=245p     
+     Cgbo=430p     Cj=720u      Cjsw=255p     Mjsw=0.3     
+     Fc=0           Tpg=-1.0
+     Theta=0.12     Eta=0.02     Kappa=10.0
*+     Wd=0.78u
*+     Rsh=150

cc4 3 1 1.1113e-14
cc11 4 0 1.8504e-13
cc49 6 7 1.2e-14
cc87 6 0 4.064e-14
cc126 11 0 9.2344e-14
cc175 7 0 2.6992e-14
cc213 14 6 1.4824e-14
cc261 4 15 3.1439e-14
cc300 17 4 1.024e-14
cc342 6 15 2.2623e-14
cc343 19 4 2.032e-14
cc344 14 0 2.6992e-14
cc345 20 0 4.6678e-14
cc383 6 17 1.2464e-14
cc384 11 15 1.288e-14
cc419 6 19 3.0648e-14
cc459 11 19 1.0982e-14
cc466 1 4 3.2832e-14
cc470 15 0 1.26282e-13
cc507 19 7 1.2e-14
cc510 17 0 4.3232e-14
cc541 1 6 1.36302e-13
cc544 19 0 4.5296e-14
cc588 11 1 2.2752e-14
cc592 3 0 1.067e-14
cc628 1 7 4.49e-14
cc668 14 19 2.1766e-14
cc672 1 0 1.79232e-13
cc675 27 28 1.65984e-13
cc760 17 15 1.024e-14
cc777 32 1 1.5288e-14
cc797 14 1 7.8984e-14
cc803 1 20 4.4738e-14
cc804 19 15 2.3232e-14
cc845 19 17 1.2688e-14
cc915 27 0 1.24008e-13
cc938 1 15 4.2789e-14
cc939 6 4 1.8768e-14
cc942 20 34 1.584e-14
cc982 1 17 3.2202e-14
cc983 11 4 1.2e-14
cc1008 37 0 1.0924e-14
cc1022 1 19 1.31805e-13
cc1049 28 0 1.16796e-13
c0 38 0 1.2301e-14
c1 1 0 3.388e-12
c2 39 0 1.2301e-14
c3 40 0 1.2301e-14
c4 41 0 1.2301e-14
c5 42 0 1.2301e-14
c6 43 0 1.2301e-14
c7 44 0 1.2301e-14
c8 45 0 1.2301e-14
c9 46 0 1.2301e-14
c10 47 0 1.2301e-14
c11 48 0 1.2301e-14
c12 49 0 1.2301e-14
c13 50 0 1.2301e-14
c14 51 0 1.2301e-14
c15 52 0 1.2301e-14
c16 53 0 1.2301e-14
c17 54 0 1.2301e-14
c18 55 0 1.2301e-14
c19 56 0 1.2301e-14
c20 57 0 1.2301e-14
c21 58 0 1.2301e-14
c22 59 0 1.2301e-14
c23 60 0 1.2301e-14
c24 27 0 3.74885e-13
c25 61 0 1.0116e-14
c26 62 0 1.2148e-14
c27 63 0 1.0116e-14
c28 64 0 1.2148e-14
c29 65 0 1.0116e-14
c30 66 0 1.2148e-14
c31 67 0 1.0116e-14
c32 68 0 1.2148e-14
c33 69 0 1.0116e-14
c34 70 0 1.2148e-14
c35 71 0 1.0116e-14
c36 72 0 1.2148e-14
c37 73 0 1.0116e-14
c38 74 0 1.2148e-14
c39 75 0 1.0116e-14
c40 76 0 1.2148e-14
c41 77 0 1.0116e-14
c42 78 0 1.2148e-14
c43 79 0 1.0116e-14
c44 80 0 1.2148e-14
c45 81 0 1.0116e-14
c46 82 0 1.2148e-14
c47 83 0 1.0116e-14
c48 84 0 1.2148e-14
c49 85 0 1.0116e-14
c50 86 0 1.2148e-14
c51 87 0 1.0116e-14
c52 88 0 1.2148e-14
c53 89 0 1.0116e-14
c54 90 0 1.2148e-14
c55 91 0 1.0116e-14
c56 92 0 1.2148e-14
c57 93 0 1.0116e-14
c58 94 0 1.2148e-14
c59 95 0 1.0116e-14
c60 96 0 1.2148e-14
c61 97 0 1.0116e-14
c62 98 0 1.2148e-14
c63 99 0 1.0116e-14
c64 100 0 1.2148e-14
c65 101 0 1.0116e-14
c66 102 0 1.2148e-14
c67 103 0 1.0116e-14
c68 104 0 1.2148e-14
c69 105 0 1.0116e-14
c70 106 0 1.2148e-14
c71 107 0 1.0116e-14
c72 108 0 1.3108e-14
c73 37 0 6.2074e-14
c74 109 0 1.1282e-14
c75 110 0 2.2644e-14
c76 111 0 8.0774e-14
c77 112 0 3.297e-14
c79 28 0 3.85102e-13
c80 113 0 3.7197e-14
c81 114 0 1.4262e-14
c82 115 0 2.7294e-14
c83 116 0 3.4903e-14
c84 117 0 3.2074e-14
c85 118 0 4.0114e-14
c86 19 0 5.55497e-13
c87 119 0 3.8458e-14
c88 120 0 1.3092e-14
c89 15 0 5.66346e-13
c91 6 0 5.6416e-13
c94 17 0 2.56302e-13
c96 14 0 2.82304e-13
c98 4 0 5.4241e-13
c103 11 0 2.63118e-13
c105 121 0 5.0108e-14
c109 122 0 2.3174e-14
c110 123 0 1.2956e-14
c111 124 0 1.5468e-14
c116 125 0 1.06678e-13
c118 7 0 1.91906e-13
c121 32 0 2.7238e-14
c123 126 0 3.4004e-14
c124 127 0 3.3074e-14
c128 128 0 2.218e-14
c132 129 0 1.2934e-14
c133 130 0 1.355e-14
c135 131 0 1.1069e-13
c138 132 0 3.6373e-14
c139 3 0 4.1085e-14
c142 133 0 1.018e-14
c144 34 0 4.2488e-14
c145 20 0 3.83758e-13
m0 1 38 149 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m1 1 39 150 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m2 1 40 151 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m3 1 41 152 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m4 1 42 153 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m5 1 43 154 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m6 1 44 155 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m7 1 45 156 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m8 1 46 157 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m9 1 47 158 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m10 1 48 159 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m11 1 49 160 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m12 1 50 161 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m13 1 51 162 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m14 1 52 163 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m15 1 53 164 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m16 1 54 165 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m17 1 55 166 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m18 1 56 167 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m19 1 57 168 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m20 1 58 169 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m21 1 59 170 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m22 1 60 171 1 pfet l=1.6e-06 w=8e-06 
+ as=4.8e-12 ad=1.4044e-10 ps=9.2e-06 pd=6.109e-05 
+ nrs=0.07 nrd=2.19 
m23 1 0 27 1 npfet l=1.6e-06 w=2.8e-06 
+ as=6.26e-12 ad=4.915e-11 ps=4.58e-06 pd=2.138e-05 
+ nrs=0.8 nrd=6.27 
m24 149 61 62 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m25 150 63 64 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m26 151 65 66 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m27 152 67 68 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m28 153 69 70 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m29 154 71 72 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m30 155 73 74 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m31 156 75 76 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m32 157 77 78 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m33 158 79 80 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m34 159 81 82 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m35 160 83 84 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m36 161 85 86 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m37 162 87 88 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m38 163 89 90 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m39 164 91 92 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m40 165 93 94 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m41 166 95 96 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m42 167 97 98 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m43 168 99 100 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m44 169 101 102 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m45 170 103 104 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m46 171 105 106 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=4.8e-12 ps=2.32e-05 pd=9.2e-06 
+ nrs=0.42 nrd=0.07 
m47 1 107 108 1 pfet l=1.6e-06 w=8e-06 
+ as=2.688e-11 ad=1.4044e-10 ps=2.32e-05 pd=6.109e-05 
+ nrs=0.42 nrd=2.19 
m48 1 37 109 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.723e-11 ad=1.1937e-10 ps=1.413e-05 pd=5.193e-05 
+ nrs=0.37 nrd=2.58 
m49 109 110 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=1.723e-11 ps=5.193e-05 pd=1.413e-05 
+ nrs=2.58 nrd=0.37 
m50 109 111 112 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.567e-11 ad=1.723e-11 ps=1.425e-05 pd=1.413e-05 
+ nrs=0.34 nrd=0.37 
m51 112 109 111 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.567e-11 ps=2.08e-05 pd=1.425e-05 
+ nrs=0.53 nrd=0.34 
m52 172 111 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.08e-05 
+ nrs=2.58 nrd=0.53 
m53 0 38 62 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m54 62 61 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m55 0 39 64 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m56 64 63 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m57 0 40 66 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m58 66 65 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m59 0 41 68 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m60 68 67 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m61 0 42 70 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m62 70 69 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m63 0 43 72 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m64 72 71 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m65 0 44 74 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m66 74 73 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m67 0 45 76 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m68 76 75 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m69 0 46 78 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m70 78 77 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m71 0 47 80 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m72 80 79 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m73 0 48 82 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m74 82 81 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m75 0 49 84 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m76 84 83 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m77 0 50 86 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m78 86 85 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m79 0 51 88 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m80 88 87 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m81 0 52 90 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m82 90 89 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m83 0 53 92 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m84 92 91 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m85 0 54 94 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m86 94 93 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m87 0 55 96 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m88 96 95 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m89 0 56 98 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m90 98 97 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m91 0 57 100 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m92 100 99 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m93 0 58 102 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m94 102 101 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m95 0 59 104 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m96 104 103 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m97 0 60 106 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.6e-12 ad=9.206e-11 ps=8.8e-06 pd=4.311e-05 
+ nrs=0.42 nrd=4 
m98 106 105 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=9.6e-12 ps=4.311e-05 pd=8.8e-06 
+ nrs=4 nrd=0.42 
m99 108 107 0 0 nfet l=1.6e-06 w=4.8e-06 
+ as=9.206e-11 ad=1.728e-11 ps=4.311e-05 pd=1.68e-05 
+ nrs=4 nrd=0.75 
m100 28 62 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m101 27 62 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m102 28 62 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m103 28 64 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m104 27 64 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m105 28 64 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m106 28 66 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m107 27 66 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m108 28 66 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m109 28 68 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m110 27 68 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m111 28 68 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m112 28 70 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m113 27 70 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m114 28 70 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m115 28 72 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m116 27 72 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m117 28 72 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m118 28 74 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m119 27 74 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m120 28 74 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m121 28 76 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m122 27 76 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m123 28 76 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m124 28 78 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m125 27 78 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m126 28 78 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m127 28 80 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m128 27 80 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m129 28 80 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m130 28 82 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m131 27 82 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m132 28 82 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m133 28 84 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m134 27 84 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m135 28 84 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m136 28 86 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m137 27 86 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m138 28 86 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m139 28 88 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m140 27 88 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m141 28 88 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m142 28 90 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m143 27 90 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m144 28 90 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m145 28 92 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m146 27 92 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m147 28 92 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m148 28 94 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m149 27 94 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m150 28 94 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m151 28 96 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m152 27 96 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m153 28 96 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m154 28 98 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m155 27 98 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m156 28 98 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m157 28 100 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m158 27 100 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m159 28 100 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m160 28 102 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m161 27 102 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m162 28 102 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m163 28 104 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m164 27 104 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m165 28 104 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m166 28 106 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m167 27 106 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m168 28 106 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m169 28 108 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m170 27 108 28 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.791e-11 ad=2.842e-11 ps=1.973e-05 pd=2.011e-05 
+ nrs=0.22 nrd=0.23 
m171 28 108 27 0 nfet l=1.6e-06 w=1.12e-05 
+ as=2.842e-11 ad=2.791e-11 ps=2.011e-05 pd=1.973e-05 
+ nrs=0.23 nrd=0.22 
m172 109 37 173 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=2.514e-11 ps=8e-06 pd=2.143e-05 
+ nrs=0.09 nrd=0.54 
m173 173 110 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=4.08e-12 ps=6.108e-05 pd=8e-06 
+ nrs=2.82 nrd=0.09 
m174 109 172 112 0 nfet l=1.6e-06 w=6.4e-06 
+ as=1.536e-11 ad=2.366e-11 ps=1.408e-05 pd=2.017e-05 
+ nrs=0.38 nrd=0.58 
m175 1 113 114 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.496e-11 ad=1.1937e-10 ps=1.12e-05 pd=5.193e-05 
+ nrs=0.32 nrd=2.58 
m176 114 115 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=1.496e-11 ps=5.193e-05 pd=1.12e-05 
+ nrs=2.58 nrd=0.32 
m177 1 114 116 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.1937e-10 ps=2.339e-05 pd=5.193e-05 
+ nrs=0.53 nrd=2.58 
m178 1 116 117 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.677e-11 ad=1.1937e-10 ps=1.457e-05 pd=5.193e-05 
+ nrs=0.36 nrd=2.58 
m179 117 118 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=1.677e-11 ps=5.193e-05 pd=1.457e-05 
+ nrs=2.58 nrd=0.36 
m180 112 109 172 0 nfet l=1.6e-06 w=6.4e-06 
+ as=2.366e-11 ad=1.536e-11 ps=2.017e-05 pd=1.408e-05 
+ nrs=0.58 nrd=0.38 
m181 172 111 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=2.514e-11 ps=6.108e-05 pd=2.143e-05 
+ nrs=2.82 nrd=0.54 
m182 114 113 174 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=2.448e-11 ps=8e-06 pd=2.08e-05 
+ nrs=0.09 nrd=0.53 
m183 120 19 119 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.152e-11 ps=1.101e-05 pd=1.36e-05 
+ nrs=1.13 nrd=1.13 
m184 116 114 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=2.448e-11 ps=6.108e-05 pd=2.339e-05 
+ nrs=2.82 nrd=0.53 
m185 117 116 175 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=2.448e-11 ps=8e-06 pd=2.339e-05 
+ nrs=0.09 nrd=0.53 
m186 174 115 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=4.08e-12 ps=6.108e-05 pd=8e-06 
+ nrs=2.82 nrd=0.09 
m187 175 118 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=4.08e-12 ps=6.108e-05 pd=8e-06 
+ nrs=2.82 nrd=0.09 
m188 120 15 119 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.152e-11 ps=1.101e-05 pd=1.36e-05 
+ nrs=1.13 nrd=1.13 
m189 0 176 111 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.3041e-10 ps=2.08e-05 pd=6.108e-05 
+ nrs=0.53 nrd=2.82 
m190 1 6 27 1 pfet l=1.6e-06 w=2e-05 
+ as=4.473e-11 ad=3.5109e-10 ps=3.27e-05 pd=0.00015273 
+ nrs=0.11 nrd=0.88 
m191 27 15 176 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.12e-12 ps=1.36e-05 pd=5.75e-06 
+ nrs=1.13 nrd=0.79 
m192 0 178 177 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.3041e-10 ps=2.339e-05 pd=6.108e-05 
+ nrs=0.53 nrd=2.82 
m193 0 111 179 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.92e-12 ad=6.137e-11 ps=4.4e-06 pd=2.874e-05 
+ nrs=0.19 nrd=5.99 
m194 179 17 180 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.92e-12 ps=9.33e-06 pd=4.4e-06 
+ nrs=0.79 nrd=0.19 
m195 0 37 180 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=6.137e-11 ps=9.33e-06 pd=2.874e-05 
+ nrs=0.79 nrd=5.99 
m196 180 14 181 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=6.4e-12 ad=8.11e-12 ps=7.2e-06 pd=9.33e-06 
+ nrs=0.63 nrd=0.79 
m197 181 4 178 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=6.4e-12 ps=1.36e-05 pd=7.2e-06 
+ nrs=1.13 nrd=0.63 
m198 27 6 1 1 pfet l=1.6e-06 w=2e-05 
+ as=3.5109e-10 ad=4.473e-11 ps=0.00015273 pd=3.27e-05 
+ nrs=0.88 nrd=0.11 
m199 27 19 176 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=7.16e-12 ps=1.36e-05 pd=5.23e-06 
+ nrs=1.13 nrd=0.7 
m200 0 183 182 0 nnfet l=1.6e-06 w=4e-06 
+ as=2.336e-11 ad=7.671e-11 ps=2.08e-05 pd=3.593e-05 
+ nrs=1.46 nrd=4.79 
m201 0 182 37 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.3041e-10 ps=2.08e-05 pd=6.108e-05 
+ nrs=0.53 nrd=2.82 
m202 177 15 183 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.152e-11 ps=1.36e-05 pd=1.101e-05 
+ nrs=1.13 nrd=1.13 
m203 0 185 184 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.1e-11 ad=1.3041e-10 ps=1.686e-05 pd=6.108e-05 
+ nrs=0.45 nrd=2.82 
m204 121 11 186 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.164e-05 
+ nrs=0.79 nrd=1.13 
m205 186 14 110 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.408e-11 ad=8.11e-12 ps=1.376e-05 pd=9.33e-06 
+ nrs=1.38 nrd=0.79 
m206 186 4 185 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m207 0 187 110 0 nfet l=1.6e-06 w=4.8e-06 
+ as=2.112e-11 ad=9.206e-11 ps=2.064e-05 pd=4.311e-05 
+ nrs=0.92 nrd=4 
m208 184 15 187 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.88e-12 ps=1.36e-05 pd=7.94e-06 
+ nrs=1.13 nrd=0.96 
m209 111 176 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.08e-05 
+ nrs=2.58 nrd=0.53 
m210 1 111 188 1 pfet l=1.6e-06 w=4.8e-06 
+ as=1.216e-11 ad=8.426e-11 ps=1.147e-05 pd=3.666e-05 
+ nrs=0.53 nrd=3.66 
m211 188 17 1 1 pfet l=1.6e-06 w=4.8e-06 
+ as=8.426e-11 ad=1.216e-11 ps=3.666e-05 pd=1.147e-05 
+ nrs=3.66 nrd=0.53 
m212 188 37 181 1 pfet l=1.6e-06 w=4.8e-06 
+ as=1.344e-11 ad=1.216e-11 ps=1.29e-05 pd=1.147e-05 
+ nrs=0.58 nrd=0.53 
m213 1 14 181 1 pfet l=1.6e-06 w=4.8e-06 
+ as=1.344e-11 ad=8.426e-11 ps=1.29e-05 pd=3.666e-05 
+ nrs=0.58 nrd=3.66 
m214 181 6 178 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.96e-12 ps=1.36e-05 pd=8.6e-06 
+ nrs=1.13 nrd=0.88 
m215 177 19 183 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.152e-11 ps=1.36e-05 pd=1.101e-05 
+ nrs=1.13 nrd=1.13 
m216 177 178 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.339e-05 
+ nrs=2.58 nrd=0.53 
m217 121 14 186 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.164e-05 
+ nrs=0.79 nrd=1.13 
m218 186 11 110 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.408e-11 ad=8.11e-12 ps=1.376e-05 pd=9.33e-06 
+ nrs=1.38 nrd=0.79 
m219 182 183 1 1 npfet l=1.6e-06 w=4e-06 
+ as=7.022e-11 ad=2.336e-11 ps=3.055e-05 pd=2.08e-05 
+ nrs=4.39 nrd=1.46 
m220 37 182 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.08e-05 
+ nrs=2.58 nrd=0.53 
m221 0 189 122 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.3041e-10 ps=2.339e-05 pd=6.108e-05 
+ nrs=0.53 nrd=2.82 
m222 124 14 123 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m223 186 6 185 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m224 184 19 187 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.88e-12 ps=1.36e-05 pd=7.94e-06 
+ nrs=1.13 nrd=0.96 
m225 184 185 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.1e-11 ps=5.193e-05 pd=1.686e-05 
+ nrs=2.58 nrd=0.45 
m226 0 191 190 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.1e-11 ad=1.3041e-10 ps=1.686e-05 pd=6.108e-05 
+ nrs=0.45 nrd=2.82 
m227 189 15 190 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=9.88e-12 ad=1.152e-11 ps=7.94e-06 pd=1.36e-05 
+ nrs=0.96 nrd=1.13 
m228 0 192 119 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.3041e-10 ps=2.339e-05 pd=6.108e-05 
+ nrs=0.53 nrd=2.82 
m229 191 4 193 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.36e-05 
+ nrs=0.79 nrd=1.13 
m230 122 14 193 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.101e-05 
+ nrs=0.79 nrd=1.13 
m231 193 11 116 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.101e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m232 0 125 194 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=6.137e-11 ps=9.33e-06 pd=2.874e-05 
+ nrs=0.79 nrd=5.99 
m233 194 7 0 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=6.137e-11 ad=8.11e-12 ps=2.874e-05 pd=9.33e-06 
+ nrs=5.99 nrd=0.79 
m234 194 120 195 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.088e-11 ad=8.11e-12 ps=1e-05 pd=9.33e-06 
+ nrs=1.06 nrd=0.79 
m235 195 14 196 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.088e-11 ps=9.33e-06 pd=1e-05 
+ nrs=0.79 nrd=1.06 
m236 196 11 117 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.101e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m237 196 4 192 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m238 124 11 123 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=8.11e-12 ps=9.33e-06 pd=9.33e-06 
+ nrs=0.79 nrd=0.79 
m239 123 14 1 1 npfet l=1.6e-06 w=3.2e-06 
+ as=5.617e-11 ad=8.11e-12 ps=2.444e-05 pd=9.33e-06 
+ nrs=5.49 nrd=0.79 
m240 110 187 1 1 pfet l=1.6e-06 w=4.8e-06 
+ as=8.426e-11 ad=2.112e-11 ps=3.666e-05 pd=2.064e-05 
+ nrs=3.66 nrd=0.92 
m241 189 19 190 1 npfet l=1.6e-06 w=3.2e-06 
+ as=9.88e-12 ad=1.152e-11 ps=7.94e-06 pd=1.36e-05 
+ nrs=0.96 nrd=1.13 
m242 122 189 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.339e-05 
+ nrs=2.58 nrd=0.53 
m243 191 6 193 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.36e-05 
+ nrs=0.79 nrd=1.13 
m244 190 191 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.1e-11 ps=5.193e-05 pd=1.686e-05 
+ nrs=2.58 nrd=0.45 
m245 122 11 193 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.101e-05 
+ nrs=0.79 nrd=1.13 
m246 193 14 116 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.101e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m247 1 125 197 1 pfet l=1.6e-06 w=5.2e-06 
+ as=3.12e-12 ad=9.128e-11 ps=6.4e-06 pd=3.971e-05 
+ nrs=0.12 nrd=3.38 
m248 197 7 195 1 pfet l=1.6e-06 w=5.2e-06 
+ as=1.236e-11 ad=3.12e-12 ps=1.224e-05 pd=6.4e-06 
+ nrs=0.46 nrd=0.12 
m249 195 120 1 1 pfet l=1.6e-06 w=5.2e-06 
+ as=9.128e-11 ad=1.236e-11 ps=3.971e-05 pd=1.224e-05 
+ nrs=3.38 nrd=0.46 
m250 1 6 28 1 pfet l=1.6e-06 w=3.36e-05 
+ as=1.2096e-10 ad=5.8983e-10 ps=7.44e-05 pd=0.00025659 
+ nrs=0.11 nrd=0.52 
m251 126 32 198 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.36e-05 
+ nrs=0.79 nrd=1.13 
m252 198 127 121 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.164e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m253 1 200 199 1 npfet l=1.6e-06 w=4e-06 
+ as=1.369e-11 ad=7.022e-11 ps=1.2e-05 pd=3.055e-05 
+ nrs=0.86 nrd=4.39 
m254 198 6 200 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m255 1 201 121 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=1.1937e-10 ps=2.473e-05 pd=5.193e-05 
+ nrs=0.53 nrd=2.58 
m256 199 19 201 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.095e-11 ps=1.36e-05 pd=9.6e-06 
+ nrs=1.13 nrd=1.07 
m257 112 7 124 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=7.38e-12 ps=9.33e-06 pd=6.7e-06 
+ nrs=0.79 nrd=0.72 
m258 124 17 128 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.12e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m259 0 15 28 0 nfet l=1.6e-06 w=8.4e-06 
+ as=2.094e-11 ad=1.611e-10 ps=1.48e-05 pd=7.545e-05 
+ nrs=0.3 nrd=2.28 
m260 28 15 0 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.611e-10 ad=2.094e-11 ps=7.545e-05 pd=1.48e-05 
+ nrs=2.28 nrd=0.3 
m261 0 15 28 0 nfet l=1.6e-06 w=8.4e-06 
+ as=2.094e-11 ad=1.611e-10 ps=1.48e-05 pd=7.545e-05 
+ nrs=0.3 nrd=2.28 
m262 28 15 0 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.611e-10 ad=2.094e-11 ps=7.545e-05 pd=1.48e-05 
+ nrs=2.28 nrd=0.3 
m263 0 15 28 0 nfet l=1.6e-06 w=8.4e-06 
+ as=2.094e-11 ad=1.611e-10 ps=1.48e-05 pd=7.545e-05 
+ nrs=0.3 nrd=2.28 
m264 28 15 0 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.611e-10 ad=2.094e-11 ps=7.545e-05 pd=1.48e-05 
+ nrs=2.28 nrd=0.3 
m265 0 15 28 0 nfet l=1.6e-06 w=8.4e-06 
+ as=2.094e-11 ad=1.611e-10 ps=1.48e-05 pd=7.545e-05 
+ nrs=0.3 nrd=2.28 
m266 28 15 0 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.611e-10 ad=2.094e-11 ps=7.545e-05 pd=1.48e-05 
+ nrs=2.28 nrd=0.3 
m267 126 127 198 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.36e-05 
+ nrs=0.79 nrd=1.13 
m268 198 32 121 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.164e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m269 198 4 200 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m270 199 15 201 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.095e-11 ps=1.36e-05 pd=9.6e-06 
+ nrs=1.13 nrd=1.07 
m271 199 200 0 0 nnfet l=1.6e-06 w=4e-06 
+ as=7.671e-11 ad=1.369e-11 ps=3.593e-05 pd=1.2e-05 
+ nrs=4.79 nrd=0.86 
m272 1 203 202 1 npfet l=1.6e-06 w=4e-06 
+ as=1.227e-11 ad=7.022e-11 ps=1.111e-05 pd=3.055e-05 
+ nrs=0.77 nrd=4.39 
m273 123 6 203 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m274 1 204 128 1 pfet l=1.6e-06 w=6.4e-06 
+ as=2.304e-11 ad=1.1235e-10 ps=2.24e-05 pd=4.887e-05 
+ nrs=0.56 nrd=2.74 
m275 1 128 129 1 pfet l=1.6e-06 w=6.4e-06 
+ as=2.304e-11 ad=1.1235e-10 ps=2e-05 pd=4.887e-05 
+ nrs=0.56 nrd=2.74 
m276 202 19 204 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.81e-12 ps=1.36e-05 pd=8.89e-06 
+ nrs=1.13 nrd=0.96 
m277 1 129 130 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.558e-11 ad=1.1937e-10 ps=1.716e-05 pd=5.193e-05 
+ nrs=0.55 nrd=2.58 
m278 130 122 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.558e-11 ps=5.193e-05 pd=1.716e-05 
+ nrs=2.58 nrd=0.55 
m279 130 7 205 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.204e-11 ps=9.33e-06 pd=8.08e-06 
+ nrs=0.79 nrd=1.18 
m280 205 17 131 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.343e-11 ad=8.11e-12 ps=1.161e-05 pd=9.33e-06 
+ nrs=1.31 nrd=0.79 
m281 112 17 124 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=7.68e-12 ps=9.33e-06 pd=7.04e-06 
+ nrs=0.79 nrd=0.75 
m282 124 7 128 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.12e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m283 123 4 203 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=1.152e-11 ps=1.36e-05 pd=1.36e-05 
+ nrs=1.13 nrd=1.13 
m284 121 201 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=2.448e-11 ps=6.108e-05 pd=2.473e-05 
+ nrs=2.82 nrd=0.53 
m285 202 15 204 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.81e-12 ps=1.36e-05 pd=8.89e-06 
+ nrs=1.13 nrd=0.96 
m286 202 203 0 0 nnfet l=1.6e-06 w=4e-06 
+ as=7.671e-11 ad=1.227e-11 ps=3.593e-05 pd=1.111e-05 
+ nrs=4.79 nrd=0.77 
m287 128 204 0 0 nfet l=1.6e-06 w=6.4e-06 
+ as=1.2274e-10 ad=2.304e-11 ps=5.748e-05 pd=2.24e-05 
+ nrs=3 nrd=0.56 
m288 129 128 0 0 nfet l=1.6e-06 w=6.4e-06 
+ as=1.2274e-10 ad=2.304e-11 ps=5.748e-05 pd=2e-05 
+ nrs=3 nrd=0.56 
m289 1 207 206 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.1e-11 ad=1.1937e-10 ps=1.686e-05 pd=5.193e-05 
+ nrs=0.45 nrd=2.58 
m290 205 6 207 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m291 195 11 196 1 npfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=7.6e-12 ps=9.33e-06 pd=7.53e-06 
+ nrs=0.79 nrd=0.74 
m292 196 14 117 1 npfet l=1.6e-06 w=3.2e-06 
+ as=7.89e-12 ad=8.11e-12 ps=6.86e-06 pd=9.33e-06 
+ nrs=0.77 nrd=0.79 
m293 196 6 192 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m294 3 119 132 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.949e-11 ad=1.949e-11 ps=1.472e-05 pd=1.472e-05 
+ nrs=0.28 nrd=0.28 
m295 132 119 3 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.949e-11 ad=1.949e-11 ps=1.472e-05 pd=1.472e-05 
+ nrs=0.28 nrd=0.28 
m296 3 119 132 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.949e-11 ad=1.949e-11 ps=1.472e-05 pd=1.472e-05 
+ nrs=0.28 nrd=0.28 
m297 132 119 3 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.949e-11 ad=1.949e-11 ps=1.472e-05 pd=1.472e-05 
+ nrs=0.28 nrd=0.28 
m298 3 119 132 0 nfet l=1.6e-06 w=8.4e-06 
+ as=1.949e-11 ad=1.949e-11 ps=1.472e-05 pd=1.472e-05 
+ nrs=0.28 nrd=0.28 
m299 119 192 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=2.448e-11 ps=5.193e-05 pd=2.339e-05 
+ nrs=2.58 nrd=0.53 
m300 131 6 208 1 npfet l=1.6e-06 w=4e-06 
+ as=2.336e-11 ad=1.678e-11 ps=2.08e-05 pd=1.451e-05 
+ nrs=1.46 nrd=1.05 
m301 1 208 209 1 pfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=1.1937e-10 ps=8e-06 pd=5.193e-05 
+ nrs=0.09 nrd=2.58 
m302 209 19 210 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=4.08e-12 ps=2.08e-05 pd=8e-06 
+ nrs=0.53 nrd=0.09 
m303 1 210 211 1 pfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=1.1937e-10 ps=8e-06 pd=5.193e-05 
+ nrs=0.09 nrd=2.58 
m304 211 6 133 1 pfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=4.08e-12 ps=2.08e-05 pd=8e-06 
+ nrs=0.53 nrd=0.09 
m305 1 133 212 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.36e-11 ad=1.1937e-10 ps=1.08e-05 pd=5.193e-05 
+ nrs=0.29 nrd=2.58 
m306 212 133 1 1 pfet l=1.6e-06 w=6.8e-06 
+ as=1.1937e-10 ad=1.36e-11 ps=5.193e-05 pd=1.08e-05 
+ nrs=2.58 nrd=0.29 
m307 1 212 34 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m308 34 212 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m309 1 34 20 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m310 20 34 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m311 1 34 20 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m312 20 34 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m313 1 34 20 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m314 20 34 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m315 1 34 20 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m316 20 34 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m317 1 34 20 1 pfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=2.8087e-10 ps=2e-05 pd=0.00012218 
+ nrs=0.13 nrd=1.1 
m318 20 34 1 1 pfet l=1.6e-06 w=1.6e-05 
+ as=2.8087e-10 ad=3.2e-11 ps=0.00012218 pd=2e-05 
+ nrs=1.1 nrd=0.13 
m319 1 213 131 1 pfet l=1.6e-06 w=1e-05 
+ as=4.195e-11 ad=1.7554e-10 ps=3.628e-05 pd=7.636e-05 
+ nrs=0.42 nrd=1.76 
m320 206 19 213 1 npfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.88e-12 ps=1.36e-05 pd=7.94e-06 
+ nrs=1.13 nrd=0.96 
m321 131 4 208 0 nnfet l=1.6e-06 w=4e-06 
+ as=2.336e-11 ad=1.678e-11 ps=2.08e-05 pd=1.451e-05 
+ nrs=1.46 nrd=1.05 
m322 0 208 214 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=1.3041e-10 ps=8e-06 pd=6.108e-05 
+ nrs=0.09 nrd=2.82 
m323 214 15 210 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=4.08e-12 ps=2.08e-05 pd=8e-06 
+ nrs=0.53 nrd=0.09 
m324 0 210 215 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=1.3041e-10 ps=8e-06 pd=6.108e-05 
+ nrs=0.09 nrd=2.82 
m325 215 4 133 0 nfet l=1.6e-06 w=6.8e-06 
+ as=2.448e-11 ad=4.08e-12 ps=2.08e-05 pd=8e-06 
+ nrs=0.53 nrd=0.09 
m326 0 133 212 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.36e-11 ad=1.3041e-10 ps=1.08e-05 pd=6.108e-05 
+ nrs=0.29 nrd=2.82 
m327 212 133 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=1.36e-11 ps=6.108e-05 pd=1.08e-05 
+ nrs=2.82 nrd=0.29 
m328 130 17 205 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=8.11e-12 ad=1.152e-11 ps=9.33e-06 pd=1.101e-05 
+ nrs=0.79 nrd=1.13 
m329 205 7 131 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.343e-11 ad=8.11e-12 ps=1.161e-05 pd=9.33e-06 
+ nrs=1.31 nrd=0.79 
m330 205 4 207 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=8.11e-12 ps=1.36e-05 pd=9.33e-06 
+ nrs=1.13 nrd=0.79 
m331 130 122 216 0 nfet l=1.6e-06 w=6.8e-06 
+ as=4.08e-12 ad=2.448e-11 ps=8e-06 pd=2.339e-05 
+ nrs=0.09 nrd=0.53 
m332 216 129 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=4.08e-12 ps=6.108e-05 pd=8e-06 
+ nrs=2.82 nrd=0.09 
m333 206 15 213 0 nnfet l=1.6e-06 w=3.2e-06 
+ as=1.152e-11 ad=9.88e-12 ps=1.36e-05 pd=7.94e-06 
+ nrs=1.13 nrd=0.96 
m334 206 207 0 0 nfet l=1.6e-06 w=6.8e-06 
+ as=1.3041e-10 ad=2.1e-11 ps=6.108e-05 pd=1.686e-05 
+ nrs=2.82 nrd=0.45 
m335 131 213 0 0 nfet l=1.6e-06 w=1e-05 
+ as=1.9179e-10 ad=4.195e-11 ps=8.982e-05 pd=3.628e-05 
+ nrs=1.92 nrd=0.42 
m336 0 212 34 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m337 34 212 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
m338 0 34 20 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m339 20 34 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
m340 0 34 20 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m341 20 34 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
m342 0 34 20 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m343 20 34 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
m344 0 34 20 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m345 20 34 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
m346 0 34 20 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.2e-11 ad=3.0686e-10 ps=2e-05 pd=0.00014371 
+ nrs=0.13 nrd=1.2 
m347 20 34 0 0 nfet l=1.6e-06 w=1.6e-05 
+ as=3.0686e-10 ad=3.2e-11 ps=0.00014371 pd=2e-05 
+ nrs=1.2 nrd=0.13 
cload 20 0 3.5e-12
VPh1H 15 0 pwl (9.3e-11 -0.003 2.36e-10 -0.005 7.85e-10 -0.022 9.28e-10 -0.026 
+ 1.131e-09 -0.019 1.274e-09 0.001 1.476e-09 0.057 1.62e-09 0.125 
+ 1.822e-09 0.274 1.966e-09 0.425 2.168e-09 0.693 2.311e-09 0.906 
+ 2.346e-09 0.96 2.37e-09 0.998 2.487e-09 1.185 2.742e-09 1.6 
+ 2.839e-09 1.758 2.977e-09 1.979 3.074e-09 2.13 3.289e-09 2.452 
+ 3.441e-09 2.667 3.657e-09 2.946 3.809e-09 3.125 4.024e-09 3.353 
+ 4.177e-09 3.494 4.392e-09 3.67 4.545e-09 3.778 4.76e-09 3.912 
+ 4.912e-09 3.993 5.128e-09 4.089 5.28e-09 4.148 5.333e-09 4.166 
+ 5.476e-09 4.211 5.55e-09 4.232 5.761e-09 4.284 5.911e-09 4.314 
+ 6.122e-09 4.35 6.271e-09 4.371 6.681e-09 4.416 6.971e-09 4.438 
+ 7.176e-09 4.449 7.322e-09 4.456 7.527e-09 4.462 8.32e-09 4.484 
+ 8.582e-09 4.501 8.767e-09 4.517 9.029e-09 4.535 9.214e-09 4.521 
+ 9.475e-09 4.455 9.66e-09 4.362 9.922e-09 4.168 1.0107e-08 3.978 
+ 1.0369e-08 3.624 1.0554e-08 3.305 1.0815e-08 2.764 1.1e-08 2.341 
+ 1.1131e-08 2.029 1.1224e-08 1.809 1.1354e-08 1.505 1.1447e-08 1.294 
+ 1.1654e-08 0.88 1.1801e-08 0.645 1.2008e-08 0.4 1.2154e-08 0.28 
+ 1.2361e-08 0.171 1.2508e-08 0.122 1.2715e-08 0.081 1.2861e-08 0.063 
+ 1.3179e-08 0.039 1.3403e-08 0.027 1.3562e-08 0.021 2.5e-08 -0.003 
+ 2.5236e-08 -0.005 2.5785e-08 -0.022 2.5928e-08 -0.026 2.6131e-08 -0.019 
+ 2.6274e-08 0.001 2.6476e-08 0.057 2.662e-08 0.125 2.6822e-08 0.274 
+ 2.6966e-08 0.425 2.7168e-08 0.693 2.7311e-08 0.906 2.7346e-08 0.96 
+ 2.737e-08 0.998 2.7487e-08 1.185 2.7742e-08 1.6 2.7839e-08 1.758 
+ 2.7977e-08 1.979 2.8074e-08 2.13 2.8289e-08 2.452 2.8441e-08 2.667 
+ 2.8657e-08 2.946 2.8809e-08 3.125 2.9024e-08 3.353 2.9177e-08 3.494 
+ 2.9392e-08 3.67 2.9545e-08 3.778 2.976e-08 3.912 2.9912e-08 3.993 
+ 3.0128e-08 4.089 3.028e-08 4.148 3.0333e-08 4.166 3.0476e-08 4.211 
+ 3.055e-08 4.232 3.0761e-08 4.284 3.0911e-08 4.314 3.1122e-08 4.35 
+ 3.1271e-08 4.371 3.1681e-08 4.416 3.1971e-08 4.438 3.2176e-08 4.449 
+ 3.2322e-08 4.456 3.2527e-08 4.462 3.332e-08 4.484 3.3582e-08 4.501 
+ 3.3767e-08 4.517 3.4029e-08 4.535 3.4214e-08 4.521 3.4475e-08 4.455 
+ 3.466e-08 4.362 3.4922e-08 4.168 3.5107e-08 3.978 3.5369e-08 3.624 
+ 3.5554e-08 3.305 3.5815e-08 2.764 3.6e-08 2.341 3.6131e-08 2.029 
+ 3.6224e-08 1.809 3.6354e-08 1.505 3.6447e-08 1.294 3.6654e-08 0.88 
+ 3.6801e-08 0.645 3.7008e-08 0.4 3.7154e-08 0.28 3.7361e-08 0.171 
+ 3.7508e-08 0.122 3.7715e-08 0.081 3.7861e-08 0.063 3.8179e-08 0.039 
+ 3.8403e-08 0.027 3.8562e-08 0.021 5e-08 -0.003 5.0236e-08 -0.005 
+ 5.0785e-08 -0.022 5.0928e-08 -0.026 5.1131e-08 -0.019 5.1274e-08 0.001 
+ 5.1476e-08 0.057 5.162e-08 0.125 5.1822e-08 0.274 5.1966e-08 0.425 
+ 5.2168e-08 0.693 5.2311e-08 0.906 5.2346e-08 0.96 5.237e-08 0.998 
+ 5.2487e-08 1.185 5.2742e-08 1.6 5.2839e-08 1.758 5.2977e-08 1.979 
+ 5.3074e-08 2.13 5.3289e-08 2.452 5.3441e-08 2.667 5.3657e-08 2.946 
+ 5.3809e-08 3.125 5.4024e-08 3.353 5.4177e-08 3.494 5.4392e-08 3.67 
+ 5.4545e-08 3.778 5.476e-08 3.912 5.4912e-08 3.993 5.5128e-08 4.089 
+ 5.528e-08 4.148 5.5333e-08 4.166 5.5476e-08 4.211 5.555e-08 4.232 
+ 5.5761e-08 4.284 5.5911e-08 4.314 5.6122e-08 4.35 5.6271e-08 4.371 
+ 5.6681e-08 4.416 5.6971e-08 4.438 5.7176e-08 4.449 5.7322e-08 4.456 
+ 5.7527e-08 4.462 5.832e-08 4.484 5.8582e-08 4.501 5.8767e-08 4.517 
+ 5.9029e-08 4.535 5.9214e-08 4.521 5.9475e-08 4.455 5.966e-08 4.362 
+ 5.9922e-08 4.168 6.0107e-08 3.978 6.0369e-08 3.624 6.0554e-08 3.305 
+ 6.0815e-08 2.764 6.1e-08 2.341 6.1131e-08 2.029 6.1224e-08 1.809 
+ 6.1354e-08 1.505 6.1447e-08 1.294 6.1654e-08 0.88 6.1801e-08 0.645 
+ 6.2008e-08 0.4 6.2154e-08 0.28 6.2361e-08 0.171 6.2508e-08 0.122 
+ 6.2715e-08 0.081 6.2861e-08 0.063 6.3179e-08 0.039 6.3403e-08 0.027 
+ 6.3562e-08 0.021 7.5e-08 -0.003 7.5236e-08 -0.005 7.5785e-08 -0.022 
+ 7.5928e-08 -0.026 7.6131e-08 -0.019 7.6274e-08 0.001 7.6476e-08 0.057 
+ 7.662e-08 0.125 7.6822e-08 0.274 7.6966e-08 0.425 7.7168e-08 0.693 
+ 7.7311e-08 0.906 7.7346e-08 0.96 7.737e-08 0.998 7.7487e-08 1.185 
+ 7.7742e-08 1.6 7.7839e-08 1.758 7.7977e-08 1.979 7.8074e-08 2.13 
+ 7.8289e-08 2.452 7.8441e-08 2.667 7.8657e-08 2.946 7.8809e-08 3.125 
+ 7.9024e-08 3.353 7.9177e-08 3.494 7.9392e-08 3.67 7.9545e-08 3.778 
+ 7.976e-08 3.912 7.9912e-08 3.993 8.0128e-08 4.089 8.028e-08 4.148 
+ 8.0333e-08 4.166 8.0476e-08 4.211 8.055e-08 4.232 8.0761e-08 4.284 
+ 8.0911e-08 4.314 8.1122e-08 4.35 8.1271e-08 4.371 8.1681e-08 4.416 
+ 8.1971e-08 4.438 8.2176e-08 4.449 8.2322e-08 4.456 8.2527e-08 4.462 
+ 8.332e-08 4.484 8.3582e-08 4.501 8.3767e-08 4.517 8.4029e-08 4.535 
+ 8.4214e-08 4.521 8.4475e-08 4.455 8.466e-08 4.362 8.4922e-08 4.168 
+ 8.5107e-08 3.978 8.5369e-08 3.624 8.5554e-08 3.305 8.5815e-08 2.764 
+ 8.6e-08 2.341 8.6131e-08 2.029 8.6224e-08 1.809 8.6354e-08 1.505 
+ 8.6447e-08 1.294 8.6654e-08 0.88 8.6801e-08 0.645 8.7008e-08 0.4 
+ 8.7154e-08 0.28 8.7361e-08 0.171 8.7508e-08 0.122 8.7715e-08 0.081 
+ 8.7861e-08 0.063 8.8179e-08 0.039 8.8403e-08 0.027 8.8562e-08 0.021 
+ 1e-07 -0.003 1.00236e-07 -0.005 1.00785e-07 -0.022 1.00928e-07 -0.026 
+ 1.01131e-07 -0.019 1.01274e-07 0.001 1.01476e-07 0.057 1.0162e-07 0.125 
+ 1.01822e-07 0.274 1.01966e-07 0.425 1.02168e-07 0.693 1.02311e-07 0.906 
+ 1.02346e-07 0.96 1.0237e-07 0.998 1.02487e-07 1.185 1.02742e-07 1.6 
+ 1.02839e-07 1.758 1.02977e-07 1.979 1.03074e-07 2.13 1.03289e-07 2.452 
+ 1.03441e-07 2.667 1.03657e-07 2.946 1.03809e-07 3.125 1.04024e-07 3.353 
+ 1.04177e-07 3.494 1.04392e-07 3.67 1.04545e-07 3.778 1.0476e-07 3.912 
+ 1.04912e-07 3.993 1.05128e-07 4.089 1.0528e-07 4.148 1.05333e-07 4.166 
+ 1.05476e-07 4.211 1.0555e-07 4.232 1.05761e-07 4.284 1.05911e-07 4.314 
+ 1.06122e-07 4.35 1.06271e-07 4.371 1.06681e-07 4.416 1.06971e-07 4.438 
+ 1.07176e-07 4.449 1.07322e-07 4.456 1.07527e-07 4.462 1.0832e-07 4.484 
+ 1.08582e-07 4.501 1.08767e-07 4.517 1.09029e-07 4.535 1.09214e-07 4.521 
+ 1.09475e-07 4.455 1.0966e-07 4.362 1.09922e-07 4.168 1.10107e-07 3.978 
+ 1.10369e-07 3.624 1.10554e-07 3.305 1.10815e-07 2.764 1.11e-07 2.341 
+ 1.11131e-07 2.029 1.11224e-07 1.809 1.11354e-07 1.505 1.11447e-07 1.294 
+ 1.11654e-07 0.88 1.11801e-07 0.645 1.12008e-07 0.4 1.12154e-07 0.28 
+ 1.12361e-07 0.171 1.12508e-07 0.122 1.12715e-07 0.081 1.12861e-07 0.063 
+ 1.13179e-07 0.039 1.13403e-07 0.027 1.13562e-07 0.021 1.25e-07 -0.003 
+ 1.25236e-07 -0.005 1.25785e-07 -0.022 1.25928e-07 -0.026 1.26131e-07 -0.019 
+ 1.26274e-07 0.001 1.26476e-07 0.057 1.2662e-07 0.125 1.26822e-07 0.274 
+ 1.26966e-07 0.425 1.27168e-07 0.693 1.27311e-07 0.906 1.27346e-07 0.96 
+ 1.2737e-07 0.998 1.27487e-07 1.185 1.27742e-07 1.6 1.27839e-07 1.758 
+ 1.27977e-07 1.979 1.28074e-07 2.13 1.28289e-07 2.452 1.28441e-07 2.667 
+ 1.28657e-07 2.946 1.28809e-07 3.125 1.29024e-07 3.353 1.29177e-07 3.494 
+ 1.29392e-07 3.67 1.29545e-07 3.778 1.2976e-07 3.912 1.29912e-07 3.993 
+ 1.30128e-07 4.089 1.3028e-07 4.148 1.30333e-07 4.166 1.30476e-07 4.211 
+ 1.3055e-07 4.232 1.30761e-07 4.284 1.30911e-07 4.314 1.31122e-07 4.35 
+ 1.31271e-07 4.371 1.31681e-07 4.416 1.31971e-07 4.438 1.32176e-07 4.449 
+ 1.32322e-07 4.456 1.32527e-07 4.462 1.3332e-07 4.484 1.33582e-07 4.501 
+ 1.33767e-07 4.517 1.34029e-07 4.535 1.34214e-07 4.521 1.34475e-07 4.455 
+ 1.3466e-07 4.362 1.34922e-07 4.168 1.35107e-07 3.978 1.35369e-07 3.624 
+ 1.35554e-07 3.305 1.35815e-07 2.764 1.36e-07 2.341 1.36131e-07 2.029 
+ 1.36224e-07 1.809 1.36354e-07 1.505 1.36447e-07 1.294 1.36654e-07 0.88 
+ 1.36801e-07 0.645 1.37008e-07 0.4 1.37154e-07 0.28 1.37361e-07 0.171 
+ 1.37508e-07 0.122 1.37715e-07 0.081 1.37861e-07 0.063 1.38179e-07 0.039 
+ 1.38403e-07 0.027 1.38562e-07 0.021 1.5e-07 -0.003 1.50236e-07 -0.005 
+ 1.50785e-07 -0.022 1.50928e-07 -0.026 1.51131e-07 -0.019 1.51274e-07 0.001 
+ 1.51476e-07 0.057 1.5162e-07 0.125 1.51822e-07 0.274 1.51966e-07 0.425 
+ 1.52168e-07 0.693 1.52311e-07 0.906 1.52346e-07 0.96 1.5237e-07 0.998 
+ 1.52487e-07 1.185 1.52742e-07 1.6 1.52839e-07 1.758 1.52977e-07 1.979 
+ 1.53074e-07 2.13 1.53289e-07 2.452 1.53441e-07 2.667 1.53657e-07 2.946 
+ 1.53809e-07 3.125 1.54024e-07 3.353 1.54177e-07 3.494 1.54392e-07 3.67 
+ 1.54545e-07 3.778 1.5476e-07 3.912 1.54912e-07 3.993 1.55128e-07 4.089 
+ 1.5528e-07 4.148 1.55333e-07 4.166 1.55476e-07 4.211 1.5555e-07 4.232 
+ 1.55761e-07 4.284 1.55911e-07 4.314 1.56122e-07 4.35 1.56271e-07 4.371 
+ 1.56681e-07 4.416 1.56971e-07 4.438 1.57176e-07 4.449 1.57322e-07 4.456 
+ 1.57527e-07 4.462 1.5832e-07 4.484 1.58582e-07 4.501 1.58767e-07 4.517 
+ 1.59029e-07 4.535 1.59214e-07 4.521 1.59475e-07 4.455 1.5966e-07 4.362 
+ 1.59922e-07 4.168 1.60107e-07 3.978 1.60369e-07 3.624 1.60554e-07 3.305 
+ 1.60815e-07 2.764 1.61e-07 2.341 1.61131e-07 2.029 1.61224e-07 1.809 
+ 1.61354e-07 1.505 1.61447e-07 1.294 1.61654e-07 0.88 1.61801e-07 0.645 
+ 1.62008e-07 0.4 1.62154e-07 0.28 1.62361e-07 0.171 1.62508e-07 0.122 
+ 1.62715e-07 0.081 1.62861e-07 0.063 1.63179e-07 0.039 1.63403e-07 0.027 
+ 1.63562e-07 0.021 1.75e-07 -0.003 1.75236e-07 -0.005 1.75785e-07 -0.022 
+ 1.75928e-07 -0.026 1.76131e-07 -0.019 1.76274e-07 0.001 1.76476e-07 0.057 
+ 1.7662e-07 0.125 1.76822e-07 0.274 1.76966e-07 0.425 1.77168e-07 0.693 
+ 1.77311e-07 0.906 1.77346e-07 0.96 1.7737e-07 0.998 1.77487e-07 1.185 
+ 1.77742e-07 1.6 1.77839e-07 1.758 1.77977e-07 1.979 1.78074e-07 2.13 
+ 1.78289e-07 2.452 1.78441e-07 2.667 1.78657e-07 2.946 1.78809e-07 3.125 
+ 1.79024e-07 3.353 1.79177e-07 3.494 1.79392e-07 3.67 1.79545e-07 3.778 
+ 1.7976e-07 3.912 1.79912e-07 3.993 1.80128e-07 4.089 1.8028e-07 4.148 
+ 1.80333e-07 4.166 1.80476e-07 4.211 1.8055e-07 4.232 1.80761e-07 4.284 
+ 1.80911e-07 4.314 1.81122e-07 4.35 1.81271e-07 4.371 1.81681e-07 4.416 
+ 1.81971e-07 4.438 1.82176e-07 4.449 1.82322e-07 4.456 1.82527e-07 4.462 
+ 1.8332e-07 4.484 1.83582e-07 4.501 1.83767e-07 4.517 1.84029e-07 4.535 
+ 1.84214e-07 4.521 1.84475e-07 4.455 1.8466e-07 4.362 1.84922e-07 4.168 
+ 1.85107e-07 3.978 1.85369e-07 3.624 1.85554e-07 3.305 1.85815e-07 2.764 
+ 1.86e-07 2.341 1.86131e-07 2.029 1.86224e-07 1.809 1.86354e-07 1.505 
+ 1.86447e-07 1.294 1.86654e-07 0.88 1.86801e-07 0.645 1.87008e-07 0.4 
+ 1.87154e-07 0.28 1.87361e-07 0.171 1.87508e-07 0.122 1.87715e-07 0.081 
+ 1.87861e-07 0.063 1.88179e-07 0.039 1.88403e-07 0.027 1.88562e-07 0.021 
+ 2e-07 -0.003 )
VPh1L 19 0 pwl (9.3e-11 4.51 2.36e-10 4.517 4.39e-10 4.528 7.85e-10 4.541 
+ 9.28e-10 4.526 1.131e-09 4.478 1.274e-09 4.421 1.476e-09 4.304 
+ 1.62e-09 4.197 1.822e-09 4.003 1.966e-09 3.833 2.168e-09 3.538 
+ 2.311e-09 3.288 2.346e-09 3.223 2.37e-09 3.176 2.439e-09 3.038 
+ 2.487e-09 2.936 2.556e-09 2.788 2.605e-09 2.68 2.742e-09 2.362 
+ 2.839e-09 2.134 3.289e-09 1.105 3.441e-09 0.82 3.657e-09 0.5 
+ 3.809e-09 0.337 4.024e-09 0.184 4.177e-09 0.117 4.392e-09 0.062 
+ 4.545e-09 0.039 4.76e-09 0.021 4.912e-09 0.014 5.128e-09 0.008 
+ 5.28e-09 0.005 8.197e-09 -0.002 8.32e-09 -0.006 8.582e-09 -0.018 
+ 8.767e-09 -0.031 9.029e-09 -0.019 9.214e-09 0.035 9.475e-09 0.2 
+ 9.66e-09 0.398 9.922e-09 0.772 1.0107e-08 1.067 1.0369e-08 1.504 
+ 1.0554e-08 1.809 1.0815e-08 2.221 1.1e-08 2.494 1.1131e-08 2.678 
+ 1.1224e-08 2.8 1.1354e-08 2.961 1.1447e-08 3.069 1.1654e-08 3.287 
+ 1.1801e-08 3.421 1.2008e-08 3.585 1.2154e-08 3.687 1.2361e-08 3.814 
+ 1.2508e-08 3.893 1.2715e-08 3.989 1.2861e-08 4.046 1.3179e-08 4.149 
+ 1.3403e-08 4.206 1.3562e-08 4.24 1.3674e-08 4.261 1.3832e-08 4.288 
+ 1.3945e-08 4.306 1.4103e-08 4.328 1.4216e-08 4.342 1.4374e-08 4.36 
+ 1.4486e-08 4.371 1.4645e-08 4.386 2.4883e-08 4.503 2.5e-08 4.51 
+ 2.5236e-08 4.517 2.5439e-08 4.528 2.5785e-08 4.541 2.5928e-08 4.526 
+ 2.6131e-08 4.478 2.6274e-08 4.421 2.6476e-08 4.304 2.662e-08 4.197 
+ 2.6822e-08 4.003 2.6966e-08 3.833 2.7168e-08 3.538 2.7311e-08 3.288 
+ 2.7346e-08 3.223 2.737e-08 3.176 2.7439e-08 3.038 2.7487e-08 2.936 
+ 2.7556e-08 2.788 2.7605e-08 2.68 2.7742e-08 2.362 2.7839e-08 2.134 
+ 2.8289e-08 1.105 2.8441e-08 0.82 2.8657e-08 0.5 2.8809e-08 0.337 
+ 2.9024e-08 0.184 2.9177e-08 0.117 2.9392e-08 0.062 2.9545e-08 0.039 
+ 2.976e-08 0.021 2.9912e-08 0.014 3.0128e-08 0.008 3.028e-08 0.005 
+ 3.3197e-08 -0.002 3.332e-08 -0.006 3.3582e-08 -0.018 3.3767e-08 -0.031 
+ 3.4029e-08 -0.019 3.4214e-08 0.035 3.4475e-08 0.2 3.466e-08 0.398 
+ 3.4922e-08 0.772 3.5107e-08 1.067 3.5369e-08 1.504 3.5554e-08 1.809 
+ 3.5815e-08 2.221 3.6e-08 2.494 3.6131e-08 2.678 3.6224e-08 2.8 
+ 3.6354e-08 2.961 3.6447e-08 3.069 3.6654e-08 3.287 3.6801e-08 3.421 
+ 3.7008e-08 3.585 3.7154e-08 3.687 3.7361e-08 3.814 3.7508e-08 3.893 
+ 3.7715e-08 3.989 3.7861e-08 4.046 3.8179e-08 4.149 3.8403e-08 4.206 
+ 3.8562e-08 4.24 3.8674e-08 4.261 3.8832e-08 4.288 3.8945e-08 4.306 
+ 3.9103e-08 4.328 3.9216e-08 4.342 3.9374e-08 4.36 3.9486e-08 4.371 
+ 3.9645e-08 4.386 4.9883e-08 4.503 5e-08 4.51 5.0236e-08 4.517 
+ 5.0439e-08 4.528 5.0785e-08 4.541 5.0928e-08 4.526 5.1131e-08 4.478 
+ 5.1274e-08 4.421 5.1476e-08 4.304 5.162e-08 4.197 5.1822e-08 4.003 
+ 5.1966e-08 3.833 5.2168e-08 3.538 5.2311e-08 3.288 5.2346e-08 3.223 
+ 5.237e-08 3.176 5.2439e-08 3.038 5.2487e-08 2.936 5.2556e-08 2.788 
+ 5.2605e-08 2.68 5.2742e-08 2.362 5.2839e-08 2.134 5.3289e-08 1.105 
+ 5.3441e-08 0.82 5.3657e-08 0.5 5.3809e-08 0.337 5.4024e-08 0.184 
+ 5.4177e-08 0.117 5.4392e-08 0.062 5.4545e-08 0.039 5.476e-08 0.021 
+ 5.4912e-08 0.014 5.5128e-08 0.008 5.528e-08 0.005 5.8197e-08 -0.002 
+ 5.832e-08 -0.006 5.8582e-08 -0.018 5.8767e-08 -0.031 5.9029e-08 -0.019 
+ 5.9214e-08 0.035 5.9475e-08 0.2 5.966e-08 0.398 5.9922e-08 0.772 
+ 6.0107e-08 1.067 6.0369e-08 1.504 6.0554e-08 1.809 6.0815e-08 2.221 
+ 6.1e-08 2.494 6.1131e-08 2.678 6.1224e-08 2.8 6.1354e-08 2.961 
+ 6.1447e-08 3.069 6.1654e-08 3.287 6.1801e-08 3.421 6.2008e-08 3.585 
+ 6.2154e-08 3.687 6.2361e-08 3.814 6.2508e-08 3.893 6.2715e-08 3.989 
+ 6.2861e-08 4.046 6.3179e-08 4.149 6.3403e-08 4.206 6.3562e-08 4.24 
+ 6.3674e-08 4.261 6.3832e-08 4.288 6.3945e-08 4.306 6.4103e-08 4.328 
+ 6.4216e-08 4.342 6.4374e-08 4.36 6.4486e-08 4.371 6.4645e-08 4.386 
+ 7.4883e-08 4.503 7.5e-08 4.51 7.5236e-08 4.517 7.5439e-08 4.528 
+ 7.5785e-08 4.541 7.5928e-08 4.526 7.6131e-08 4.478 7.6274e-08 4.421 
+ 7.6476e-08 4.304 7.662e-08 4.197 7.6822e-08 4.003 7.6966e-08 3.833 
+ 7.7168e-08 3.538 7.7311e-08 3.288 7.7346e-08 3.223 7.737e-08 3.176 
+ 7.7439e-08 3.038 7.7487e-08 2.936 7.7556e-08 2.788 7.7605e-08 2.68 
+ 7.7742e-08 2.362 7.7839e-08 2.134 7.8289e-08 1.105 7.8441e-08 0.82 
+ 7.8657e-08 0.5 7.8809e-08 0.337 7.9024e-08 0.184 7.9177e-08 0.117 
+ 7.9392e-08 0.062 7.9545e-08 0.039 7.976e-08 0.021 7.9912e-08 0.014 
+ 8.0128e-08 0.008 8.028e-08 0.005 8.3197e-08 -0.002 8.332e-08 -0.006 
+ 8.3582e-08 -0.018 8.3767e-08 -0.031 8.4029e-08 -0.019 8.4214e-08 0.035 
+ 8.4475e-08 0.2 8.466e-08 0.398 8.4922e-08 0.772 8.5107e-08 1.067 
+ 8.5369e-08 1.504 8.5554e-08 1.809 8.5815e-08 2.221 8.6e-08 2.494 
+ 8.6131e-08 2.678 8.6224e-08 2.8 8.6354e-08 2.961 8.6447e-08 3.069 
+ 8.6654e-08 3.287 8.6801e-08 3.421 8.7008e-08 3.585 8.7154e-08 3.687 
+ 8.7361e-08 3.814 8.7508e-08 3.893 8.7715e-08 3.989 8.7861e-08 4.046 
+ 8.8179e-08 4.149 8.8403e-08 4.206 8.8562e-08 4.24 8.8674e-08 4.261 
+ 8.8832e-08 4.288 8.8945e-08 4.306 8.9103e-08 4.328 8.9216e-08 4.342 
+ 8.9374e-08 4.36 8.9486e-08 4.371 8.9645e-08 4.386 9.9883e-08 4.503 
+ 1e-07 4.51 1.00236e-07 4.517 1.00439e-07 4.528 1.00785e-07 4.541 
+ 1.00928e-07 4.526 1.01131e-07 4.478 1.01274e-07 4.421 1.01476e-07 4.304 
+ 1.0162e-07 4.197 1.01822e-07 4.003 1.01966e-07 3.833 1.02168e-07 3.538 
+ 1.02311e-07 3.288 1.02346e-07 3.223 1.0237e-07 3.176 1.02439e-07 3.038 
+ 1.02487e-07 2.936 1.02556e-07 2.788 1.02605e-07 2.68 1.02742e-07 2.362 
+ 1.02839e-07 2.134 1.03289e-07 1.105 1.03441e-07 0.82 1.03657e-07 0.5 
+ 1.03809e-07 0.337 1.04024e-07 0.184 1.04177e-07 0.117 1.04392e-07 0.062 
+ 1.04545e-07 0.039 1.0476e-07 0.021 1.04912e-07 0.014 1.05128e-07 0.008 
+ 1.0528e-07 0.005 1.08197e-07 -0.002 1.0832e-07 -0.006 1.08582e-07 -0.018 
+ 1.08767e-07 -0.031 1.09029e-07 -0.019 1.09214e-07 0.035 1.09475e-07 0.2 
+ 1.0966e-07 0.398 1.09922e-07 0.772 1.10107e-07 1.067 1.10369e-07 1.504 
+ 1.10554e-07 1.809 1.10815e-07 2.221 1.11e-07 2.494 1.11131e-07 2.678 
+ 1.11224e-07 2.8 1.11354e-07 2.961 1.11447e-07 3.069 1.11654e-07 3.287 
+ 1.11801e-07 3.421 1.12008e-07 3.585 1.12154e-07 3.687 1.12361e-07 3.814 
+ 1.12508e-07 3.893 1.12715e-07 3.989 1.12861e-07 4.046 1.13179e-07 4.149 
+ 1.13403e-07 4.206 1.13562e-07 4.24 1.13674e-07 4.261 1.13832e-07 4.288 
+ 1.13945e-07 4.306 1.14103e-07 4.328 1.14216e-07 4.342 1.14374e-07 4.36 
+ 1.14486e-07 4.371 1.14645e-07 4.386 1.24883e-07 4.503 1.25e-07 4.51 
+ 1.25236e-07 4.517 1.25439e-07 4.528 1.25785e-07 4.541 1.25928e-07 4.526 
+ 1.26131e-07 4.478 1.26274e-07 4.421 1.26476e-07 4.304 1.2662e-07 4.197 
+ 1.26822e-07 4.003 1.26966e-07 3.833 1.27168e-07 3.538 1.27311e-07 3.288 
+ 1.27346e-07 3.223 1.2737e-07 3.176 1.27439e-07 3.038 1.27487e-07 2.936 
+ 1.27556e-07 2.788 1.27605e-07 2.68 1.27742e-07 2.362 1.27839e-07 2.134 
+ 1.28289e-07 1.105 1.28441e-07 0.82 1.28657e-07 0.5 1.28809e-07 0.337 
+ 1.29024e-07 0.184 1.29177e-07 0.117 1.29392e-07 0.062 1.29545e-07 0.039 
+ 1.2976e-07 0.021 1.29912e-07 0.014 1.30128e-07 0.008 1.3028e-07 0.005 
+ 1.33197e-07 -0.002 1.3332e-07 -0.006 1.33582e-07 -0.018 1.33767e-07 -0.031 
+ 1.34029e-07 -0.019 1.34214e-07 0.035 1.34475e-07 0.2 1.3466e-07 0.398 
+ 1.34922e-07 0.772 1.35107e-07 1.067 1.35369e-07 1.504 1.35554e-07 1.809 
+ 1.35815e-07 2.221 1.36e-07 2.494 1.36131e-07 2.678 1.36224e-07 2.8 
+ 1.36354e-07 2.961 1.36447e-07 3.069 1.36654e-07 3.287 1.36801e-07 3.421 
+ 1.37008e-07 3.585 1.37154e-07 3.687 1.37361e-07 3.814 1.37508e-07 3.893 
+ 1.37715e-07 3.989 1.37861e-07 4.046 1.38179e-07 4.149 1.38403e-07 4.206 
+ 1.38562e-07 4.24 1.38674e-07 4.261 1.38832e-07 4.288 1.38945e-07 4.306 
+ 1.39103e-07 4.328 1.39216e-07 4.342 1.39374e-07 4.36 1.39486e-07 4.371 
+ 1.39645e-07 4.386 1.49883e-07 4.503 1.5e-07 4.51 1.50236e-07 4.517 
+ 1.50439e-07 4.528 1.50785e-07 4.541 1.50928e-07 4.526 1.51131e-07 4.478 
+ 1.51274e-07 4.421 1.51476e-07 4.304 1.5162e-07 4.197 1.51822e-07 4.003 
+ 1.51966e-07 3.833 1.52168e-07 3.538 1.52311e-07 3.288 1.52346e-07 3.223 
+ 1.5237e-07 3.176 1.52439e-07 3.038 1.52487e-07 2.936 1.52556e-07 2.788 
+ 1.52605e-07 2.68 1.52742e-07 2.362 1.52839e-07 2.134 1.53289e-07 1.105 
+ 1.53441e-07 0.82 1.53657e-07 0.5 1.53809e-07 0.337 1.54024e-07 0.184 
+ 1.54177e-07 0.117 1.54392e-07 0.062 1.54545e-07 0.039 1.5476e-07 0.021 
+ 1.54912e-07 0.014 1.55128e-07 0.008 1.5528e-07 0.005 1.58197e-07 -0.002 
+ 1.5832e-07 -0.006 1.58582e-07 -0.018 1.58767e-07 -0.031 1.59029e-07 -0.019 
+ 1.59214e-07 0.035 1.59475e-07 0.2 1.5966e-07 0.398 1.59922e-07 0.772 
+ 1.60107e-07 1.067 1.60369e-07 1.504 1.60554e-07 1.809 1.60815e-07 2.221 
+ 1.61e-07 2.494 1.61131e-07 2.678 1.61224e-07 2.8 1.61354e-07 2.961 
+ 1.61447e-07 3.069 1.61654e-07 3.287 1.61801e-07 3.421 1.62008e-07 3.585 
+ 1.62154e-07 3.687 1.62361e-07 3.814 1.62508e-07 3.893 1.62715e-07 3.989 
+ 1.62861e-07 4.046 1.63179e-07 4.149 1.63403e-07 4.206 1.63562e-07 4.24 
+ 1.63674e-07 4.261 1.63832e-07 4.288 1.63945e-07 4.306 1.64103e-07 4.328 
+ 1.64216e-07 4.342 1.64374e-07 4.36 1.64486e-07 4.371 1.64645e-07 4.386 
+ 1.74883e-07 4.503 1.75e-07 4.51 1.75236e-07 4.517 1.75439e-07 4.528 
+ 1.75785e-07 4.541 1.75928e-07 4.526 1.76131e-07 4.478 1.76274e-07 4.421 
+ 1.76476e-07 4.304 1.7662e-07 4.197 1.76822e-07 4.003 1.76966e-07 3.833 
+ 1.77168e-07 3.538 1.77311e-07 3.288 1.77346e-07 3.223 1.7737e-07 3.176 
+ 1.77439e-07 3.038 1.77487e-07 2.936 1.77556e-07 2.788 1.77605e-07 2.68 
+ 1.77742e-07 2.362 1.77839e-07 2.134 1.78289e-07 1.105 1.78441e-07 0.82 
+ 1.78657e-07 0.5 1.78809e-07 0.337 1.79024e-07 0.184 1.79177e-07 0.117 
+ 1.79392e-07 0.062 1.79545e-07 0.039 1.7976e-07 0.021 1.79912e-07 0.014 
+ 1.80128e-07 0.008 1.8028e-07 0.005 1.83197e-07 -0.002 1.8332e-07 -0.006 
+ 1.83582e-07 -0.018 1.83767e-07 -0.031 1.84029e-07 -0.019 1.84214e-07 0.035 
+ 1.84475e-07 0.2 1.8466e-07 0.398 1.84922e-07 0.772 1.85107e-07 1.067 
+ 1.85369e-07 1.504 1.85554e-07 1.809 1.85815e-07 2.221 1.86e-07 2.494 
+ 1.86131e-07 2.678 1.86224e-07 2.8 1.86354e-07 2.961 1.86447e-07 3.069 
+ 1.86654e-07 3.287 1.86801e-07 3.421 1.87008e-07 3.585 1.87154e-07 3.687 
+ 1.87361e-07 3.814 1.87508e-07 3.893 1.87715e-07 3.989 1.87861e-07 4.046 
+ 1.88179e-07 4.149 1.88403e-07 4.206 1.88562e-07 4.24 1.88674e-07 4.261 
+ 1.88832e-07 4.288 1.88945e-07 4.306 1.89103e-07 4.328 1.89216e-07 4.342 
+ 1.89374e-07 4.36 1.89486e-07 4.371 1.89645e-07 4.386 1.99883e-07 4.503 
+ 2e-07 4.51 )
VPh2H 4 0 pwl (9.3e-11 0.057 2.36e-10 0.045 4.39e-10 0.033 5.82e-10 0.026 
+ 7.85e-10 0.018 1.3562e-08 -0.015 1.3674e-08 -0.021 1.3832e-08 -0.026 
+ 1.3945e-08 -0.024 1.4103e-08 -0.011 1.4216e-08 0.008 1.4374e-08 0.054 
+ 1.4486e-08 0.103 1.4645e-08 0.202 1.4757e-08 0.301 1.4823e-08 0.37 
+ 1.487e-08 0.424 1.5002e-08 0.593 1.5095e-08 0.726 1.5228e-08 0.925 
+ 1.5321e-08 1.072 1.5453e-08 1.284 1.5546e-08 1.436 1.5772e-08 1.803 
+ 1.5997e-08 2.16 1.6129e-08 2.358 1.6223e-08 2.494 1.6355e-08 2.679 
+ 1.6448e-08 2.803 1.658e-08 2.968 1.6674e-08 3.079 1.6789e-08 3.208 
+ 1.687e-08 3.294 1.71e-08 3.511 1.7263e-08 3.645 1.7493e-08 3.808 
+ 1.7655e-08 3.908 1.8011e-08 4.082 1.8263e-08 4.177 1.8619e-08 4.275 
+ 1.8871e-08 4.327 1.9227e-08 4.379 1.9479e-08 4.406 1.9657e-08 4.42 
+ 1.9783e-08 4.429 2.0087e-08 4.446 2.0719e-08 4.484 2.087e-08 4.498 
+ 2.1235e-08 4.527 2.1448e-08 4.511 2.16e-08 4.474 2.1813e-08 4.38 
+ 2.1964e-08 4.282 2.2178e-08 4.101 2.2329e-08 3.936 2.2543e-08 3.644 
+ 2.2694e-08 3.391 2.2908e-08 2.97 2.3059e-08 2.637 2.3273e-08 2.135 
+ 2.3637e-08 1.288 2.3788e-08 0.984 2.4002e-08 0.632 2.4153e-08 0.447 
+ 2.4367e-08 0.268 2.4518e-08 0.185 2.4732e-08 0.115 2.4883e-08 0.084 
+ 2.5e-08 0.057 2.5236e-08 0.045 2.5439e-08 0.033 2.5582e-08 0.026 
+ 2.5785e-08 0.018 3.8562e-08 -0.015 3.8674e-08 -0.021 3.8832e-08 -0.026 
+ 3.8945e-08 -0.024 3.9103e-08 -0.011 3.9216e-08 0.008 3.9374e-08 0.054 
+ 3.9486e-08 0.103 3.9645e-08 0.202 3.9757e-08 0.301 3.9823e-08 0.37 
+ 3.987e-08 0.424 4.0002e-08 0.593 4.0095e-08 0.726 4.0228e-08 0.925 
+ 4.0321e-08 1.072 4.0453e-08 1.284 4.0546e-08 1.436 4.0772e-08 1.803 
+ 4.0997e-08 2.16 4.1129e-08 2.358 4.1223e-08 2.494 4.1355e-08 2.679 
+ 4.1448e-08 2.803 4.158e-08 2.968 4.1674e-08 3.079 4.1789e-08 3.208 
+ 4.187e-08 3.294 4.21e-08 3.511 4.2263e-08 3.645 4.2493e-08 3.808 
+ 4.2655e-08 3.908 4.3011e-08 4.082 4.3263e-08 4.177 4.3619e-08 4.275 
+ 4.3871e-08 4.327 4.4227e-08 4.379 4.4479e-08 4.406 4.4657e-08 4.42 
+ 4.4783e-08 4.429 4.5087e-08 4.446 4.5719e-08 4.484 4.587e-08 4.498 
+ 4.6235e-08 4.527 4.6448e-08 4.511 4.66e-08 4.474 4.6813e-08 4.38 
+ 4.6964e-08 4.282 4.7178e-08 4.101 4.7329e-08 3.936 4.7543e-08 3.644 
+ 4.7694e-08 3.391 4.7908e-08 2.97 4.8059e-08 2.637 4.8273e-08 2.135 
+ 4.8637e-08 1.288 4.8788e-08 0.984 4.9002e-08 0.632 4.9153e-08 0.447 
+ 4.9367e-08 0.268 4.9518e-08 0.185 4.9732e-08 0.115 4.9883e-08 0.084 
+ 5e-08 0.057 5.0236e-08 0.045 5.0439e-08 0.033 5.0582e-08 0.026 
+ 5.0785e-08 0.018 6.3562e-08 -0.015 6.3674e-08 -0.021 6.3832e-08 -0.026 
+ 6.3945e-08 -0.024 6.4103e-08 -0.011 6.4216e-08 0.008 6.4374e-08 0.054 
+ 6.4486e-08 0.103 6.4645e-08 0.202 6.4757e-08 0.301 6.4823e-08 0.37 
+ 6.487e-08 0.424 6.5002e-08 0.593 6.5095e-08 0.726 6.5228e-08 0.925 
+ 6.5321e-08 1.072 6.5453e-08 1.284 6.5546e-08 1.436 6.5772e-08 1.803 
+ 6.5997e-08 2.16 6.6129e-08 2.358 6.6223e-08 2.494 6.6355e-08 2.679 
+ 6.6448e-08 2.803 6.658e-08 2.968 6.6674e-08 3.079 6.6789e-08 3.208 
+ 6.687e-08 3.294 6.71e-08 3.511 6.7263e-08 3.645 6.7493e-08 3.808 
+ 6.7655e-08 3.908 6.8011e-08 4.082 6.8263e-08 4.177 6.8619e-08 4.275 
+ 6.8871e-08 4.327 6.9227e-08 4.379 6.9479e-08 4.406 6.9657e-08 4.42 
+ 6.9783e-08 4.429 7.0087e-08 4.446 7.0719e-08 4.484 7.087e-08 4.498 
+ 7.1235e-08 4.527 7.1448e-08 4.511 7.16e-08 4.474 7.1813e-08 4.38 
+ 7.1964e-08 4.282 7.2178e-08 4.101 7.2329e-08 3.936 7.2543e-08 3.644 
+ 7.2694e-08 3.391 7.2908e-08 2.97 7.3059e-08 2.637 7.3273e-08 2.135 
+ 7.3637e-08 1.288 7.3788e-08 0.984 7.4002e-08 0.632 7.4153e-08 0.447 
+ 7.4367e-08 0.268 7.4518e-08 0.185 7.4732e-08 0.115 7.4883e-08 0.084 
+ 7.5e-08 0.057 7.5236e-08 0.045 7.5439e-08 0.033 7.5582e-08 0.026 
+ 7.5785e-08 0.018 8.8562e-08 -0.015 8.8674e-08 -0.021 8.8832e-08 -0.026 
+ 8.8945e-08 -0.024 8.9103e-08 -0.011 8.9216e-08 0.008 8.9374e-08 0.054 
+ 8.9486e-08 0.103 8.9645e-08 0.202 8.9757e-08 0.301 8.9823e-08 0.37 
+ 8.987e-08 0.424 9.0002e-08 0.593 9.0095e-08 0.726 9.0228e-08 0.925 
+ 9.0321e-08 1.072 9.0453e-08 1.284 9.0546e-08 1.436 9.0772e-08 1.803 
+ 9.0997e-08 2.16 9.1129e-08 2.358 9.1223e-08 2.494 9.1355e-08 2.679 
+ 9.1448e-08 2.803 9.158e-08 2.968 9.1674e-08 3.079 9.1789e-08 3.208 
+ 9.187e-08 3.294 9.21e-08 3.511 9.2263e-08 3.645 9.2493e-08 3.808 
+ 9.2655e-08 3.908 9.3011e-08 4.082 9.3263e-08 4.177 9.3619e-08 4.275 
+ 9.3871e-08 4.327 9.4227e-08 4.379 9.4479e-08 4.406 9.4657e-08 4.42 
+ 9.4783e-08 4.429 9.5087e-08 4.446 9.5719e-08 4.484 9.587e-08 4.498 
+ 9.6235e-08 4.527 9.6448e-08 4.511 9.66e-08 4.474 9.6813e-08 4.38 
+ 9.6964e-08 4.282 9.7178e-08 4.101 9.7329e-08 3.936 9.7543e-08 3.644 
+ 9.7694e-08 3.391 9.7908e-08 2.97 9.8059e-08 2.637 9.8273e-08 2.135 
+ 9.8637e-08 1.288 9.8788e-08 0.984 9.9002e-08 0.632 9.9153e-08 0.447 
+ 9.9367e-08 0.268 9.9518e-08 0.185 9.9732e-08 0.115 9.9883e-08 0.084 
+ 1e-07 0.057 1.00236e-07 0.045 1.00439e-07 0.033 1.00582e-07 0.026 
+ 1.00785e-07 0.018 1.13562e-07 -0.015 1.13674e-07 -0.021 1.13832e-07 -0.026 
+ 1.13945e-07 -0.024 1.14103e-07 -0.011 1.14216e-07 0.008 1.14374e-07 0.054 
+ 1.14486e-07 0.103 1.14645e-07 0.202 1.14757e-07 0.301 1.14823e-07 0.37 
+ 1.1487e-07 0.424 1.15002e-07 0.593 1.15095e-07 0.726 1.15228e-07 0.925 
+ 1.15321e-07 1.072 1.15453e-07 1.284 1.15546e-07 1.436 1.15772e-07 1.803 
+ 1.15997e-07 2.16 1.16129e-07 2.358 1.16223e-07 2.494 1.16355e-07 2.679 
+ 1.16448e-07 2.803 1.1658e-07 2.968 1.16674e-07 3.079 1.16789e-07 3.208 
+ 1.1687e-07 3.294 1.171e-07 3.511 1.17263e-07 3.645 1.17493e-07 3.808 
+ 1.17655e-07 3.908 1.18011e-07 4.082 1.18263e-07 4.177 1.18619e-07 4.275 
+ 1.18871e-07 4.327 1.19227e-07 4.379 1.19479e-07 4.406 1.19657e-07 4.42 
+ 1.19783e-07 4.429 1.20087e-07 4.446 1.20719e-07 4.484 1.2087e-07 4.498 
+ 1.21235e-07 4.527 1.21448e-07 4.511 1.216e-07 4.474 1.21813e-07 4.38 
+ 1.21964e-07 4.282 1.22178e-07 4.101 1.22329e-07 3.936 1.22543e-07 3.644 
+ 1.22694e-07 3.391 1.22908e-07 2.97 1.23059e-07 2.637 1.23273e-07 2.135 
+ 1.23637e-07 1.288 1.23788e-07 0.984 1.24002e-07 0.632 1.24153e-07 0.447 
+ 1.24367e-07 0.268 1.24518e-07 0.185 1.24732e-07 0.115 1.24883e-07 0.084 
+ 1.25e-07 0.057 1.25236e-07 0.045 1.25439e-07 0.033 1.25582e-07 0.026 
+ 1.25785e-07 0.018 1.38562e-07 -0.015 1.38674e-07 -0.021 1.38832e-07 -0.026 
+ 1.38945e-07 -0.024 1.39103e-07 -0.011 1.39216e-07 0.008 1.39374e-07 0.054 
+ 1.39486e-07 0.103 1.39645e-07 0.202 1.39757e-07 0.301 1.39823e-07 0.37 
+ 1.3987e-07 0.424 1.40002e-07 0.593 1.40095e-07 0.726 1.40228e-07 0.925 
+ 1.40321e-07 1.072 1.40453e-07 1.284 1.40546e-07 1.436 1.40772e-07 1.803 
+ 1.40997e-07 2.16 1.41129e-07 2.358 1.41223e-07 2.494 1.41355e-07 2.679 
+ 1.41448e-07 2.803 1.4158e-07 2.968 1.41674e-07 3.079 1.41789e-07 3.208 
+ 1.4187e-07 3.294 1.421e-07 3.511 1.42263e-07 3.645 1.42493e-07 3.808 
+ 1.42655e-07 3.908 1.43011e-07 4.082 1.43263e-07 4.177 1.43619e-07 4.275 
+ 1.43871e-07 4.327 1.44227e-07 4.379 1.44479e-07 4.406 1.44657e-07 4.42 
+ 1.44783e-07 4.429 1.45087e-07 4.446 1.45719e-07 4.484 1.4587e-07 4.498 
+ 1.46235e-07 4.527 1.46448e-07 4.511 1.466e-07 4.474 1.46813e-07 4.38 
+ 1.46964e-07 4.282 1.47178e-07 4.101 1.47329e-07 3.936 1.47543e-07 3.644 
+ 1.47694e-07 3.391 1.47908e-07 2.97 1.48059e-07 2.637 1.48273e-07 2.135 
+ 1.48637e-07 1.288 1.48788e-07 0.984 1.49002e-07 0.632 1.49153e-07 0.447 
+ 1.49367e-07 0.268 1.49518e-07 0.185 1.49732e-07 0.115 1.49883e-07 0.084 
+ 1.5e-07 0.057 1.50236e-07 0.045 1.50439e-07 0.033 1.50582e-07 0.026 
+ 1.50785e-07 0.018 1.63562e-07 -0.015 1.63674e-07 -0.021 1.63832e-07 -0.026 
+ 1.63945e-07 -0.024 1.64103e-07 -0.011 1.64216e-07 0.008 1.64374e-07 0.054 
+ 1.64486e-07 0.103 1.64645e-07 0.202 1.64757e-07 0.301 1.64823e-07 0.37 
+ 1.6487e-07 0.424 1.65002e-07 0.593 1.65095e-07 0.726 1.65228e-07 0.925 
+ 1.65321e-07 1.072 1.65453e-07 1.284 1.65546e-07 1.436 1.65772e-07 1.803 
+ 1.65997e-07 2.16 1.66129e-07 2.358 1.66223e-07 2.494 1.66355e-07 2.679 
+ 1.66448e-07 2.803 1.6658e-07 2.968 1.66674e-07 3.079 1.66789e-07 3.208 
+ 1.6687e-07 3.294 1.671e-07 3.511 1.67263e-07 3.645 1.67493e-07 3.808 
+ 1.67655e-07 3.908 1.68011e-07 4.082 1.68263e-07 4.177 1.68619e-07 4.275 
+ 1.68871e-07 4.327 1.69227e-07 4.379 1.69479e-07 4.406 1.69657e-07 4.42 
+ 1.69783e-07 4.429 1.70087e-07 4.446 1.70719e-07 4.484 1.7087e-07 4.498 
+ 1.71235e-07 4.527 1.71448e-07 4.511 1.716e-07 4.474 1.71813e-07 4.38 
+ 1.71964e-07 4.282 1.72178e-07 4.101 1.72329e-07 3.936 1.72543e-07 3.644 
+ 1.72694e-07 3.391 1.72908e-07 2.97 1.73059e-07 2.637 1.73273e-07 2.135 
+ 1.73637e-07 1.288 1.73788e-07 0.984 1.74002e-07 0.632 1.74153e-07 0.447 
+ 1.74367e-07 0.268 1.74518e-07 0.185 1.74732e-07 0.115 1.74883e-07 0.084 
+ 1.75e-07 0.057 1.75236e-07 0.045 1.75439e-07 0.033 1.75582e-07 0.026 
+ 1.75785e-07 0.018 1.88562e-07 -0.015 1.88674e-07 -0.021 1.88832e-07 -0.026 
+ 1.88945e-07 -0.024 1.89103e-07 -0.011 1.89216e-07 0.008 1.89374e-07 0.054 
+ 1.89486e-07 0.103 1.89645e-07 0.202 1.89757e-07 0.301 1.89823e-07 0.37 
+ 1.8987e-07 0.424 1.90002e-07 0.593 1.90095e-07 0.726 1.90228e-07 0.925 
+ 1.90321e-07 1.072 1.90453e-07 1.284 1.90546e-07 1.436 1.90772e-07 1.803 
+ 1.90997e-07 2.16 1.91129e-07 2.358 1.91223e-07 2.494 1.91355e-07 2.679 
+ 1.91448e-07 2.803 1.9158e-07 2.968 1.91674e-07 3.079 1.91789e-07 3.208 
+ 1.9187e-07 3.294 1.921e-07 3.511 1.92263e-07 3.645 1.92493e-07 3.808 
+ 1.92655e-07 3.908 1.93011e-07 4.082 1.93263e-07 4.177 1.93619e-07 4.275 
+ 1.93871e-07 4.327 1.94227e-07 4.379 1.94479e-07 4.406 1.94657e-07 4.42 
+ 1.94783e-07 4.429 1.95087e-07 4.446 1.95719e-07 4.484 1.9587e-07 4.498 
+ 1.96235e-07 4.527 1.96448e-07 4.511 1.966e-07 4.474 1.96813e-07 4.38 
+ 1.96964e-07 4.282 1.97178e-07 4.101 1.97329e-07 3.936 1.97543e-07 3.644 
+ 1.97694e-07 3.391 1.97908e-07 2.97 1.98059e-07 2.637 1.98273e-07 2.135 
+ 1.98637e-07 1.288 1.98788e-07 0.984 1.99002e-07 0.632 1.99153e-07 0.447 
+ 1.99367e-07 0.268 1.99518e-07 0.185 1.99732e-07 0.115 1.99883e-07 0.084 
+ 2e-07 0.057 )
VPh2L 6 0 pwl (9.3e-11 4.116 2.36e-10 4.157 4.39e-10 4.208 5.82e-10 4.238 
+ 7.85e-10 4.275 9.28e-10 4.298 1.131e-09 4.326 1.274e-09 4.344 
+ 1.476e-09 4.366 1.62e-09 4.38 1.822e-09 4.397 1.966e-09 4.407 
+ 1.2861e-08 4.506 1.3179e-08 4.52 1.3403e-08 4.533 1.3674e-08 4.54 
+ 1.3832e-08 4.524 1.3945e-08 4.5 1.4103e-08 4.447 1.4216e-08 4.393 
+ 1.4374e-08 4.295 1.4486e-08 4.211 1.4645e-08 4.067 1.4757e-08 3.946 
+ 1.4823e-08 3.867 1.487e-08 3.806 1.5002e-08 3.617 1.5095e-08 3.466 
+ 1.5228e-08 3.227 1.5321e-08 3.041 1.5453e-08 2.759 1.5546e-08 2.548 
+ 1.5678e-08 2.238 1.5904e-08 1.706 1.5997e-08 1.489 1.6129e-08 1.191 
+ 1.6223e-08 1 1.6355e-08 0.761 1.6448e-08 0.615 1.658e-08 0.444 
+ 1.6674e-08 0.348 1.6789e-08 0.255 1.687e-08 0.203 1.71e-08 0.104 
+ 1.7263e-08 0.063 1.7493e-08 0.032 1.7655e-08 0.02 1.8011e-08 0.007 
+ 1.8263e-08 0.003 1.8619e-08 0.002 2.0332e-08 -0.005 2.0505e-08 -0.011 
+ 2.0719e-08 -0.026 2.087e-08 -0.032 2.1084e-08 -0.018 2.1235e-08 0.023 
+ 2.1448e-08 0.137 2.16e-08 0.273 2.1813e-08 0.539 2.1964e-08 0.764 
+ 2.2178e-08 1.11 2.2329e-08 1.362 2.2694e-08 1.964 2.2908e-08 2.294 
+ 2.3059e-08 2.515 2.3273e-08 2.806 2.3424e-08 2.993 2.3637e-08 3.229 
+ 2.3788e-08 3.375 2.4002e-08 3.553 2.4153e-08 3.662 2.4367e-08 3.795 
+ 2.4518e-08 3.878 2.4732e-08 3.979 2.4883e-08 4.04 2.5e-08 4.116 
+ 2.5236e-08 4.157 2.5439e-08 4.208 2.5582e-08 4.238 2.5785e-08 4.275 
+ 2.5928e-08 4.298 2.6131e-08 4.326 2.6274e-08 4.344 2.6476e-08 4.366 
+ 2.662e-08 4.38 2.6822e-08 4.397 2.6966e-08 4.407 3.7861e-08 4.506 
+ 3.8179e-08 4.52 3.8403e-08 4.533 3.8674e-08 4.54 3.8832e-08 4.524 
+ 3.8945e-08 4.5 3.9103e-08 4.447 3.9216e-08 4.393 3.9374e-08 4.295 
+ 3.9486e-08 4.211 3.9645e-08 4.067 3.9757e-08 3.946 3.9823e-08 3.867 
+ 3.987e-08 3.806 4.0002e-08 3.617 4.0095e-08 3.466 4.0228e-08 3.227 
+ 4.0321e-08 3.041 4.0453e-08 2.759 4.0546e-08 2.548 4.0678e-08 2.238 
+ 4.0904e-08 1.706 4.0997e-08 1.489 4.1129e-08 1.191 4.1223e-08 1 
+ 4.1355e-08 0.761 4.1448e-08 0.615 4.158e-08 0.444 4.1674e-08 0.348 
+ 4.1789e-08 0.255 4.187e-08 0.203 4.21e-08 0.104 4.2263e-08 0.063 
+ 4.2493e-08 0.032 4.2655e-08 0.02 4.3011e-08 0.007 4.3263e-08 0.003 
+ 4.3619e-08 0.002 4.5332e-08 -0.005 4.5505e-08 -0.011 4.5719e-08 -0.026 
+ 4.587e-08 -0.032 4.6084e-08 -0.018 4.6235e-08 0.023 4.6448e-08 0.137 
+ 4.66e-08 0.273 4.6813e-08 0.539 4.6964e-08 0.764 4.7178e-08 1.11 
+ 4.7329e-08 1.362 4.7694e-08 1.964 4.7908e-08 2.294 4.8059e-08 2.515 
+ 4.8273e-08 2.806 4.8424e-08 2.993 4.8637e-08 3.229 4.8788e-08 3.375 
+ 4.9002e-08 3.553 4.9153e-08 3.662 4.9367e-08 3.795 4.9518e-08 3.878 
+ 4.9732e-08 3.979 4.9883e-08 4.04 5e-08 4.116 5.0236e-08 4.157 
+ 5.0439e-08 4.208 5.0582e-08 4.238 5.0785e-08 4.275 5.0928e-08 4.298 
+ 5.1131e-08 4.326 5.1274e-08 4.344 5.1476e-08 4.366 5.162e-08 4.38 
+ 5.1822e-08 4.397 5.1966e-08 4.407 6.2861e-08 4.506 6.3179e-08 4.52 
+ 6.3403e-08 4.533 6.3674e-08 4.54 6.3832e-08 4.524 6.3945e-08 4.5 
+ 6.4103e-08 4.447 6.4216e-08 4.393 6.4374e-08 4.295 6.4486e-08 4.211 
+ 6.4645e-08 4.067 6.4757e-08 3.946 6.4823e-08 3.867 6.487e-08 3.806 
+ 6.5002e-08 3.617 6.5095e-08 3.466 6.5228e-08 3.227 6.5321e-08 3.041 
+ 6.5453e-08 2.759 6.5546e-08 2.548 6.5678e-08 2.238 6.5904e-08 1.706 
+ 6.5997e-08 1.489 6.6129e-08 1.191 6.6223e-08 1 6.6355e-08 0.761 
+ 6.6448e-08 0.615 6.658e-08 0.444 6.6674e-08 0.348 6.6789e-08 0.255 
+ 6.687e-08 0.203 6.71e-08 0.104 6.7263e-08 0.063 6.7493e-08 0.032 
+ 6.7655e-08 0.02 6.8011e-08 0.007 6.8263e-08 0.003 6.8619e-08 0.002 
+ 7.0332e-08 -0.005 7.0505e-08 -0.011 7.0719e-08 -0.026 7.087e-08 -0.032 
+ 7.1084e-08 -0.018 7.1235e-08 0.023 7.1448e-08 0.137 7.16e-08 0.273 
+ 7.1813e-08 0.539 7.1964e-08 0.764 7.2178e-08 1.11 7.2329e-08 1.362 
+ 7.2694e-08 1.964 7.2908e-08 2.294 7.3059e-08 2.515 7.3273e-08 2.806 
+ 7.3424e-08 2.993 7.3637e-08 3.229 7.3788e-08 3.375 7.4002e-08 3.553 
+ 7.4153e-08 3.662 7.4367e-08 3.795 7.4518e-08 3.878 7.4732e-08 3.979 
+ 7.4883e-08 4.04 7.5e-08 4.116 7.5236e-08 4.157 7.5439e-08 4.208 
+ 7.5582e-08 4.238 7.5785e-08 4.275 7.5928e-08 4.298 7.6131e-08 4.326 
+ 7.6274e-08 4.344 7.6476e-08 4.366 7.662e-08 4.38 7.6822e-08 4.397 
+ 7.6966e-08 4.407 8.7861e-08 4.506 8.8179e-08 4.52 8.8403e-08 4.533 
+ 8.8674e-08 4.54 8.8832e-08 4.524 8.8945e-08 4.5 8.9103e-08 4.447 
+ 8.9216e-08 4.393 8.9374e-08 4.295 8.9486e-08 4.211 8.9645e-08 4.067 
+ 8.9757e-08 3.946 8.9823e-08 3.867 8.987e-08 3.806 9.0002e-08 3.617 
+ 9.0095e-08 3.466 9.0228e-08 3.227 9.0321e-08 3.041 9.0453e-08 2.759 
+ 9.0546e-08 2.548 9.0678e-08 2.238 9.0904e-08 1.706 9.0997e-08 1.489 
+ 9.1129e-08 1.191 9.1223e-08 1 9.1355e-08 0.761 9.1448e-08 0.615 
+ 9.158e-08 0.444 9.1674e-08 0.348 9.1789e-08 0.255 9.187e-08 0.203 
+ 9.21e-08 0.104 9.2263e-08 0.063 9.2493e-08 0.032 9.2655e-08 0.02 
+ 9.3011e-08 0.007 9.3263e-08 0.003 9.3619e-08 0.002 9.5332e-08 -0.005 
+ 9.5505e-08 -0.011 9.5719e-08 -0.026 9.587e-08 -0.032 9.6084e-08 -0.018 
+ 9.6235e-08 0.023 9.6448e-08 0.137 9.66e-08 0.273 9.6813e-08 0.539 
+ 9.6964e-08 0.764 9.7178e-08 1.11 9.7329e-08 1.362 9.7694e-08 1.964 
+ 9.7908e-08 2.294 9.8059e-08 2.515 9.8273e-08 2.806 9.8424e-08 2.993 
+ 9.8637e-08 3.229 9.8788e-08 3.375 9.9002e-08 3.553 9.9153e-08 3.662 
+ 9.9367e-08 3.795 9.9518e-08 3.878 9.9732e-08 3.979 9.9883e-08 4.04 
+ 1e-07 4.116 1.00236e-07 4.157 1.00439e-07 4.208 1.00582e-07 4.238 
+ 1.00785e-07 4.275 1.00928e-07 4.298 1.01131e-07 4.326 1.01274e-07 4.344 
+ 1.01476e-07 4.366 1.0162e-07 4.38 1.01822e-07 4.397 1.01966e-07 4.407 
+ 1.12861e-07 4.506 1.13179e-07 4.52 1.13403e-07 4.533 1.13674e-07 4.54 
+ 1.13832e-07 4.524 1.13945e-07 4.5 1.14103e-07 4.447 1.14216e-07 4.393 
+ 1.14374e-07 4.295 1.14486e-07 4.211 1.14645e-07 4.067 1.14757e-07 3.946 
+ 1.14823e-07 3.867 1.1487e-07 3.806 1.15002e-07 3.617 1.15095e-07 3.466 
+ 1.15228e-07 3.227 1.15321e-07 3.041 1.15453e-07 2.759 1.15546e-07 2.548 
+ 1.15678e-07 2.238 1.15904e-07 1.706 1.15997e-07 1.489 1.16129e-07 1.191 
+ 1.16223e-07 1 1.16355e-07 0.761 1.16448e-07 0.615 1.1658e-07 0.444 
+ 1.16674e-07 0.348 1.16789e-07 0.255 1.1687e-07 0.203 1.171e-07 0.104 
+ 1.17263e-07 0.063 1.17493e-07 0.032 1.17655e-07 0.02 1.18011e-07 0.007 
+ 1.18263e-07 0.003 1.18619e-07 0.002 1.20332e-07 -0.005 1.20505e-07 -0.011 
+ 1.20719e-07 -0.026 1.2087e-07 -0.032 1.21084e-07 -0.018 1.21235e-07 0.023 
+ 1.21448e-07 0.137 1.216e-07 0.273 1.21813e-07 0.539 1.21964e-07 0.764 
+ 1.22178e-07 1.11 1.22329e-07 1.362 1.22694e-07 1.964 1.22908e-07 2.294 
+ 1.23059e-07 2.515 1.23273e-07 2.806 1.23424e-07 2.993 1.23637e-07 3.229 
+ 1.23788e-07 3.375 1.24002e-07 3.553 1.24153e-07 3.662 1.24367e-07 3.795 
+ 1.24518e-07 3.878 1.24732e-07 3.979 1.24883e-07 4.04 1.25e-07 4.116 
+ 1.25236e-07 4.157 1.25439e-07 4.208 1.25582e-07 4.238 1.25785e-07 4.275 
+ 1.25928e-07 4.298 1.26131e-07 4.326 1.26274e-07 4.344 1.26476e-07 4.366 
+ 1.2662e-07 4.38 1.26822e-07 4.397 1.26966e-07 4.407 1.37861e-07 4.506 
+ 1.38179e-07 4.52 1.38403e-07 4.533 1.38674e-07 4.54 1.38832e-07 4.524 
+ 1.38945e-07 4.5 1.39103e-07 4.447 1.39216e-07 4.393 1.39374e-07 4.295 
+ 1.39486e-07 4.211 1.39645e-07 4.067 1.39757e-07 3.946 1.39823e-07 3.867 
+ 1.3987e-07 3.806 1.40002e-07 3.617 1.40095e-07 3.466 1.40228e-07 3.227 
+ 1.40321e-07 3.041 1.40453e-07 2.759 1.40546e-07 2.548 1.40678e-07 2.238 
+ 1.40904e-07 1.706 1.40997e-07 1.489 1.41129e-07 1.191 1.41223e-07 1 
+ 1.41355e-07 0.761 1.41448e-07 0.615 1.4158e-07 0.444 1.41674e-07 0.348 
+ 1.41789e-07 0.255 1.4187e-07 0.203 1.421e-07 0.104 1.42263e-07 0.063 
+ 1.42493e-07 0.032 1.42655e-07 0.02 1.43011e-07 0.007 1.43263e-07 0.003 
+ 1.43619e-07 0.002 1.45332e-07 -0.005 1.45505e-07 -0.011 1.45719e-07 -0.026 
+ 1.4587e-07 -0.032 1.46084e-07 -0.018 1.46235e-07 0.023 1.46448e-07 0.137 
+ 1.466e-07 0.273 1.46813e-07 0.539 1.46964e-07 0.764 1.47178e-07 1.11 
+ 1.47329e-07 1.362 1.47694e-07 1.964 1.47908e-07 2.294 1.48059e-07 2.515 
+ 1.48273e-07 2.806 1.48424e-07 2.993 1.48637e-07 3.229 1.48788e-07 3.375 
+ 1.49002e-07 3.553 1.49153e-07 3.662 1.49367e-07 3.795 1.49518e-07 3.878 
+ 1.49732e-07 3.979 1.49883e-07 4.04 1.5e-07 4.116 1.50236e-07 4.157 
+ 1.50439e-07 4.208 1.50582e-07 4.238 1.50785e-07 4.275 1.50928e-07 4.298 
+ 1.51131e-07 4.326 1.51274e-07 4.344 1.51476e-07 4.366 1.5162e-07 4.38 
+ 1.51822e-07 4.397 1.51966e-07 4.407 1.62861e-07 4.506 1.63179e-07 4.52 
+ 1.63403e-07 4.533 1.63674e-07 4.54 1.63832e-07 4.524 1.63945e-07 4.5 
+ 1.64103e-07 4.447 1.64216e-07 4.393 1.64374e-07 4.295 1.64486e-07 4.211 
+ 1.64645e-07 4.067 1.64757e-07 3.946 1.64823e-07 3.867 1.6487e-07 3.806 
+ 1.65002e-07 3.617 1.65095e-07 3.466 1.65228e-07 3.227 1.65321e-07 3.041 
+ 1.65453e-07 2.759 1.65546e-07 2.548 1.65678e-07 2.238 1.65904e-07 1.706 
+ 1.65997e-07 1.489 1.66129e-07 1.191 1.66223e-07 1 1.66355e-07 0.761 
+ 1.66448e-07 0.615 1.6658e-07 0.444 1.66674e-07 0.348 1.66789e-07 0.255 
+ 1.6687e-07 0.203 1.671e-07 0.104 1.67263e-07 0.063 1.67493e-07 0.032 
+ 1.67655e-07 0.02 1.68011e-07 0.007 1.68263e-07 0.003 1.68619e-07 0.002 
+ 1.70332e-07 -0.005 1.70505e-07 -0.011 1.70719e-07 -0.026 1.7087e-07 -0.032 
+ 1.71084e-07 -0.018 1.71235e-07 0.023 1.71448e-07 0.137 1.716e-07 0.273 
+ 1.71813e-07 0.539 1.71964e-07 0.764 1.72178e-07 1.11 1.72329e-07 1.362 
+ 1.72694e-07 1.964 1.72908e-07 2.294 1.73059e-07 2.515 1.73273e-07 2.806 
+ 1.73424e-07 2.993 1.73637e-07 3.229 1.73788e-07 3.375 1.74002e-07 3.553 
+ 1.74153e-07 3.662 1.74367e-07 3.795 1.74518e-07 3.878 1.74732e-07 3.979 
+ 1.74883e-07 4.04 1.75e-07 4.116 1.75236e-07 4.157 1.75439e-07 4.208 
+ 1.75582e-07 4.238 1.75785e-07 4.275 1.75928e-07 4.298 1.76131e-07 4.326 
+ 1.76274e-07 4.344 1.76476e-07 4.366 1.7662e-07 4.38 1.76822e-07 4.397 
+ 1.76966e-07 4.407 1.87861e-07 4.506 1.88179e-07 4.52 1.88403e-07 4.533 
+ 1.88674e-07 4.54 1.88832e-07 4.524 1.88945e-07 4.5 1.89103e-07 4.447 
+ 1.89216e-07 4.393 1.89374e-07 4.295 1.89486e-07 4.211 1.89645e-07 4.067 
+ 1.89757e-07 3.946 1.89823e-07 3.867 1.8987e-07 3.806 1.90002e-07 3.617 
+ 1.90095e-07 3.466 1.90228e-07 3.227 1.90321e-07 3.041 1.90453e-07 2.759 
+ 1.90546e-07 2.548 1.90678e-07 2.238 1.90904e-07 1.706 1.90997e-07 1.489 
+ 1.91129e-07 1.191 1.91223e-07 1 1.91355e-07 0.761 1.91448e-07 0.615 
+ 1.9158e-07 0.444 1.91674e-07 0.348 1.91789e-07 0.255 1.9187e-07 0.203 
+ 1.921e-07 0.104 1.92263e-07 0.063 1.92493e-07 0.032 1.92655e-07 0.02 
+ 1.93011e-07 0.007 1.93263e-07 0.003 1.93619e-07 0.002 1.95332e-07 -0.005 
+ 1.95505e-07 -0.011 1.95719e-07 -0.026 1.9587e-07 -0.032 1.96084e-07 -0.018 
+ 1.96235e-07 0.023 1.96448e-07 0.137 1.966e-07 0.273 1.96813e-07 0.539 
+ 1.96964e-07 0.764 1.97178e-07 1.11 1.97329e-07 1.362 1.97694e-07 1.964 
+ 1.97908e-07 2.294 1.98059e-07 2.515 1.98273e-07 2.806 1.98424e-07 2.993 
+ 1.98637e-07 3.229 1.98788e-07 3.375 1.99002e-07 3.553 1.99153e-07 3.662 
+ 1.99367e-07 3.795 1.99518e-07 3.878 1.99732e-07 3.979 1.99883e-07 4.04 
+ 2e-07 4.116 )
VWordHSP2 127 0 pwl (0 4.5 3.75e-08 4.5 3.85e-08 0 1.875e-07 0 
+ 1.885e-07 4.5 2.125e-07 4.5 2.135e-07 0 )
VWordLSP2 32 0 pwl (0 0 3.75e-08 0 3.85e-08 4.5 1.875e-07 4.5 
+ 1.885e-07 0 2.125e-07 0 2.135e-07 4.5 )
VPostCHSP2 11 0 pwl (0 0 3.75e-08 0 4.55e-08 4.5 6.25e-08 4.5 
+ 6.75e-08 0 1.875e-07 0 2.125e-07 0 )
VPostCLSP2 14 0 pwl (0 4.5 3.75e-08 4.5 4.25e-08 0 6.25e-08 0 
+ 7.05e-08 4.5 1.875e-07 4.5 2.125e-07 4.5 )
VShiftHSP2 17 0 pwl (0 4.5 1.875e-07 4.5 3.625e-07 4.5 )
VShiftLSP2 7 0 pwl (0 0 1.875e-07 0 3.625e-07 0 )
VD31HSP2 126 0 pwl (0 4.5 3.75e-08 4.5 3.85e-08 0 1.875e-07 0 
+ 1.885e-07 4.5 2.125e-07 4.5 2.135e-07 0 )
VMBIHSP2 118 0 pwl (0 0 3.75e-08 0 3.85e-08 4.5 6.25e-08 4.5 
+ 6.35e-08 0 1.875e-07 0 2.125e-07 0 )
VABEnHSP2 113 0 pwl (0 0 3.75e-08 0 3.85e-08 4.5 6.25e-08 4.5 
+ 6.35e-08 0 1.875e-07 0 2.125e-07 0 )
VTok64LSP2 115 0 pwl (0 4.5 1.875e-07 4.5 3.625e-07 4.5 )
VTokOutLSP2 125 0 pwl (0 4.5 1.375e-07 4.5 1.385e-07 0 1.625e-07 0 
+ 1.635e-07 4.5 1.875e-07 4.5 3.125e-07 4.5 )
VMan22LSP1 39 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan21LSP1 40 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan20LSP1 41 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan19LSP1 42 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan18LSP1 43 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan17LSP1 44 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan16LSP1 45 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 1.75e-07 4.5 
+ 1.76e-07 0 2e-07 0 )
VMan15LSP1 46 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan14LSP1 47 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan13LSP1 48 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan12LSP1 49 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan11LSP1 50 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan10LSP1 51 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan9LSP1 52 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan8LSP1 53 0 pwl (0 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan7LSP1 54 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan6LSP1 55 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan5LSP1 56 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 2e-07 0 )
VMan4LSP1 57 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan3LSP1 58 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan2LSP1 59 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan1LSP1 60 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VMan0LSP1 38 0 pwl (0 0 1e-07 0 1.01e-07 4.5 1.25e-07 4.5 
+ 1.26e-07 0 1.5e-07 0 1.51e-07 4.5 2e-07 4.5 
+ 2.01e-07 0 )
VTok23LSP1 107 0 pwl (0 4.5 2e-07 4.5 )
VTok22LSP1 63 0 pwl (0 4.5 2e-07 4.5 )
VTok21LSP1 65 0 pwl (0 4.5 2e-07 4.5 )
VTok20LSP1 67 0 pwl (0 4.5 2e-07 4.5 )
VTok19LSP1 69 0 pwl (0 4.5 2e-07 4.5 )
VTok18LSP1 71 0 pwl (0 4.5 2e-07 4.5 )
VTok17LSP1 73 0 pwl (0 4.5 2e-07 4.5 )
VTok16LSP1 75 0 pwl (0 4.5 2e-07 4.5 )
VTok15LSP1 77 0 pwl (0 4.5 2e-07 4.5 )
VTok14LSP1 79 0 pwl (0 4.5 2e-07 4.5 )
VTok13LSP1 81 0 pwl (0 4.5 2e-07 4.5 )
VTok12LSP1 83 0 pwl (0 4.5 2e-07 4.5 )
VTok11LSP1 85 0 pwl (0 4.5 2e-07 4.5 )
VTok10LSP1 87 0 pwl (0 4.5 2e-07 4.5 )
VTok9LSP1 89 0 pwl (0 4.5 2e-07 4.5 )
VTok8LSP1 91 0 pwl (0 4.5 1e-07 4.5 1.01e-07 0 1.25e-07 0 
+ 1.26e-07 4.5 2e-07 4.5 )
VTok7LSP1 93 0 pwl (0 4.5 1.25e-07 4.5 1.26e-07 0 1.5e-07 0 
+ 1.51e-07 4.5 2e-07 4.5 )
VTok6LSP1 95 0 pwl (0 4.5 1.5e-07 4.5 1.51e-07 0 1.75e-07 0 
+ 1.76e-07 4.5 2e-07 4.5 )
VTok5LSP1 97 0 pwl (0 4.5 1.75e-07 4.5 1.76e-07 0 2e-07 0 
+ 2.01e-07 4.5 )
VTok4LSP1 99 0 pwl (0 4.5 2e-07 4.5 )
VTok3LSP1 101 0 pwl (0 4.5 2e-07 4.5 )
VTok2LSP1 103 0 pwl (0 4.5 2e-07 4.5 )
VTok1LSP1 105 0 pwl (0 4.5 2e-07 4.5 )
VTok0LSP1 61 0 pwl (0 4.5 2e-07 4.5 )
VVdd 1 0 4.5 
.temp 100 
.NODESET v(27)=4.5 v(28)=4.5 v(176)=4.5 v(111)=0 v(177)=4.5 v(119)=0 v(109)=0 
*.print TRAN v(15) v(4) v(127) v(11) v(17) v(28) 
+v(27) v(176) v(111) v(37) v(109) v(119) 
+v(112) v(128) v(130) v(131) v(20) 
.options limpts=50000 itl5=50000
*.TRAN 1e-09 2e-07
.end
