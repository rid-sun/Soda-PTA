mux8.sp SPICE FILE
.model nenh nmos  level = 2    vto = 0.779   kp = 3.52e-05   gamma = 1.04    phi = 0.6     cgso = 5.2e-10   cgdo = 5.2e-10    rsh = 25   cj = 0.00042    mj = 0.5   cjsw = 9e-10   mjsw = 0.33    tox = 5e-08   nsub = 1e+16    nss = 0   nfs = 1.306e+11   tpg = 1    xj = 3.85e-08   ld = 1e-07   uo = 400    ucrit = 999000   uexp = 0.001001    vmax = 32585.3   neff = 0.01001     delta = 1.33
.model penh pmos  level = 2    vto = -0.988   kp = 1.206e-05   gamma = 0.619    phi = 0.6     cgso = 4e-10   cgdo = 4e-10    rsh = 95   cj = 0.00032    mj = 0.5   cjsw = 5.5e-10   mjsw = 0.33    tox = 5e-08   nsub = 8.158e+14    nss = 0   nfs = 5.55e+09   tpg = -1    xj = 1.46e-07   ld = 2.52e-07   uo = 150    ucrit = 54941   uexp = 0.17    vmax = 100000   neff = 0.01001     delta = 1.129
m1 445 330 334 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m2 445 3314 334 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m3 335 3314 445 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m4 335 330 445 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m5 0 331 3314 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m6 1 331 3314 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m7 3314 331 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m8 1 442 331 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m9 3314 331 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m10 0 442 331 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m11 0 332 444 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m12 1 332 444 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m13 444 332 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m14 1 445 332 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m15 444 332 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m16 0 445 332 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m17 0 333 336 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m18 1 333 336 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m19 336 333 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m20 1 441 333 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m21 336 333 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m22 0 441 333 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m23 0 336 3315 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m24 1 336 3315 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m25 3315 336 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m26 3315 336 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m27 334 336 3310 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m28 334 3315 3310 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m29 3311 3315 334 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m30 3311 336 334 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m31 335 336 3312 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m32 335 3315 3312 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m33 3313 3315 335 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m34 3313 336 335 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m35 0 339 338 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m36 1 339 338 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m37 338 339 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m38 1 440 339 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m39 338 339 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m40 0 440 339 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m41 0 338 337 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m42 1 338 337 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m43 337 338 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m44 337 338 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m45 3310 338 221 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m46 3310 337 221 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m47 225 337 3310 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m48 225 338 3310 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m49 3311 338 223 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m50 3311 337 223 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m51 227 337 3311 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m52 227 338 3311 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m53 3312 338 220 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m54 3312 337 220 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m55 224 337 3312 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m56 224 338 3312 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m57 3313 338 222 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m58 3313 337 222 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
md1 226 337 3313 1 penh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m59 226 338 3313 0 nenh l=3e-06 w=7e-06   as=5.6e-11 ad=5.6e-11 ps=3e-05 pd=3e-05 
m60 330 3314 0 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m61 330 3314 1 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m62 1 3314 330 1 penh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
m63 0 3314 330 0 nenh l=3e-06 w=1.4e-05   as=1.12e-10 ad=1.12e-10 ps=4.4e-05 pd=4.4e-05 
c442 442 0 6.42e-14
c441 441 0 1.29e-13
c440 440 0 9.6e-15
c444 444 0 1.47e-14
cf1 221 0 2.259e-13
cf2 222 0 1.638e-13
cf3 223 0 2.067e-13
cf4 224 0 1.698e-13
cf5 225 0 2.127e-13
cf6 226 0 1.506e-13
cf7 227 0 1.935e-13
cf0 220 0 1.83e-13
c445 445 0 4.28e-14
c330 330 0 4.67e-14
c331 331 0 2.37e-14
c332 332 0 2.37e-14
c333 333 0 2.37e-14
c334 334 0 9.18e-14
c335 335 0 8.73e-14
c336 336 0 1.007e-13
c337 337 0 1.25e-13
c338 338 0 1.586e-13
c339 339 0 2.37e-14
c3310 3310 0 1.359e-13
c3311 3311 0 1.335e-13
c3312 3312 0 1.185e-13
c3313 3313 0 1.161e-13
c3314 3314 0 7.87e-14
c3315 3315 0 7.07e-14
vVdd 1 0 5 
V220 220 0 pwl (0 5 2e-06 5 2.001e-06 0 1.6e-05 0   1.6001e-05 5 1.8e-05 5 1.8001e-05 0 2e-05 0   2.0001e-05 5 2.2e-05 5 2.2001e-05 0 3.6e-05 0   3.6001e-05 5 3.8e-05 5 3.8001e-05 0 4e-05 0   4.0001e-05 5 4.2e-05 5 )
V221 221 0 pwl (0 0 2e-06 0 2.001e-06 5 4e-06 5   4.001e-06 0 1.8e-05 0 1.8001e-05 5 2e-05 5   2.0001e-05 0 2.2e-05 0 2.2001e-05 5 2.4e-05 5   2.4001e-05 0 3.8e-05 0 3.8001e-05 5 4e-05 5   4.0001e-05 0 4.2e-05 0 )
V222 222 0 pwl (0 0 4e-06 0 4.001e-06 5 6e-06 5   6.001e-06 0 2e-05 0 2.4e-05 0 2.4001e-05 5   2.6e-05 5 2.6001e-05 0 4e-05 0 )
V223 223 0 pwl (0 0 6e-06 0 6.001e-06 5 8e-06 5   8.001e-06 0 2e-05 0 2.6e-05 0 2.6001e-05 5   2.8e-05 5 2.8001e-05 0 4e-05 0 )
V224 224 0 pwl (0 0 8e-06 0 8.001e-06 5 1e-05 5   1.0001e-05 0 2e-05 0 2.8e-05 0 2.8001e-05 5   3e-05 5 3.0001e-05 0 4e-05 0 )
V225 225 0 pwl (0 0 1e-05 0 1.0001e-05 5 1.2e-05 5   1.2001e-05 0 2e-05 0 3e-05 0 3.0001e-05 5   3.2e-05 5 3.2001e-05 0 4e-05 0 )
V226 226 0 pwl (0 0 1.2e-05 0 1.2001e-05 5 1.4e-05 5   1.4001e-05 0 2e-05 0 3.2e-05 0 3.2001e-05 5   3.4e-05 5 3.4001e-05 0 4e-05 0 )
V227 227 0 pwl (0 0 1.4e-05 0 1.4001e-05 5 1.6e-05 5   1.6001e-05 0 2e-05 0 3.4e-05 0 3.4001e-05 5   3.6e-05 5 3.6001e-05 0 4e-05 0 )
V440 440 0 pwl (0 0 2.5e-07 0 2.51e-07 5 5e-07 5   5.01e-07 0 7.5e-07 0 7.51e-07 5 1e-06 5   1.001e-06 0 1.25e-06 0 1.251e-06 5 1.5e-06 5   1.501e-06 0 1.75e-06 0 1.751e-06 5 2e-06 5   2.001e-06 0 2.25e-06 0 2.251e-06 5 2.5e-06 5   2.501e-06 0 2.75e-06 0 2.751e-06 5 3e-06 5   3.001e-06 0 3.25e-06 0 3.251e-06 5 3.5e-06 5   3.501e-06 0 3.75e-06 0 3.751e-06 5 4e-06 5   4.001e-06 0 4.25e-06 0 4.251e-06 5 4.5e-06 5   4.501e-06 0 4.75e-06 0 4.751e-06 5 5e-06 5   5.001e-06 0 5.25e-06 0 5.251e-06 5 5.5e-06 5   5.501e-06 0 5.75e-06 0 5.751e-06 5 6e-06 5   6.001e-06 0 6.25e-06 0 6.251e-06 5 6.5e-06 5   6.501e-06 0 6.75e-06 0 6.751e-06 5 7e-06 5   7.001e-06 0 7.25e-06 0 7.251e-06 5 7.5e-06 5   7.501e-06 0 7.75e-06 0 7.751e-06 5 8e-06 5   8.001e-06 0 8.25e-06 0 8.251e-06 5 8.5e-06 5   8.501e-06 0 8.75e-06 0 8.751e-06 5 9e-06 5   9.001e-06 0 9.25e-06 0 9.251e-06 5 9.5e-06 5   9.501e-06 0 9.75e-06 0 9.751e-06 5 1e-05 5   1.0001e-05 0 1.025e-05 0 1.0251e-05 5 1.05e-05 5   1.0501e-05 0 1.075e-05 0 1.0751e-05 5 1.1e-05 5   1.1001e-05 0 1.125e-05 0 1.1251e-05 5 1.15e-05 5   1.1501e-05 0 1.175e-05 0 1.1751e-05 5 1.2e-05 5   1.2001e-05 0 1.225e-05 0 1.2251e-05 5 1.25e-05 5   1.2501e-05 0 1.275e-05 0 1.2751e-05 5 1.3e-05 5   1.3001e-05 0 1.325e-05 0 1.3251e-05 5 1.35e-05 5   1.3501e-05 0 1.375e-05 0 1.3751e-05 5 1.4e-05 5   1.4001e-05 0 1.425e-05 0 1.4251e-05 5 1.45e-05 5   1.4501e-05 0 1.475e-05 0 1.4751e-05 5 1.5e-05 5   1.5001e-05 0 1.525e-05 0 1.5251e-05 5 1.55e-05 5   1.5501e-05 0 1.575e-05 0 1.5751e-05 5 1.6e-05 5   1.6001e-05 0 1.625e-05 0 1.6251e-05 5 1.65e-05 5   1.6501e-05 0 1.675e-05 0 1.6751e-05 5 1.7e-05 5   1.7001e-05 0 1.725e-05 0 1.7251e-05 5 1.75e-05 5   1.7501e-05 0 1.775e-05 0 1.7751e-05 5 1.8e-05 5   1.8001e-05 0 1.825e-05 0 1.8251e-05 5 1.85e-05 5   1.8501e-05 0 1.875e-05 0 1.8751e-05 5 1.9e-05 5   1.9001e-05 0 1.925e-05 0 1.9251e-05 5 1.95e-05 5   1.9501e-05 0 1.975e-05 0 1.9751e-05 5 2e-05 5   2.0001e-05 0 2.025e-05 0 2.0251e-05 5 2.05e-05 5   2.0501e-05 0 2.075e-05 0 2.0751e-05 5 2.1e-05 5   2.1001e-05 0 2.125e-05 0 2.1251e-05 5 2.15e-05 5   2.1501e-05 0 2.175e-05 0 2.1751e-05 5 2.2e-05 5   2.2001e-05 0 2.225e-05 0 2.2251e-05 5 2.25e-05 5   2.2501e-05 0 2.275e-05 0 2.2751e-05 5 2.3e-05 5   2.3001e-05 0 2.325e-05 0 2.3251e-05 5 2.35e-05 5   2.3501e-05 0 2.375e-05 0 2.3751e-05 5 2.4e-05 5   2.4001e-05 0 2.425e-05 0 2.4251e-05 5 2.45e-05 5   2.4501e-05 0 2.475e-05 0 2.4751e-05 5 2.5e-05 5   2.5001e-05 0 2.525e-05 0 2.5251e-05 5 2.55e-05 5   2.5501e-05 0 2.575e-05 0 2.5751e-05 5 2.6e-05 5   2.6001e-05 0 2.625e-05 0 2.6251e-05 5 2.65e-05 5   2.6501e-05 0 2.675e-05 0 2.6751e-05 5 2.7e-05 5   2.7001e-05 0 2.725e-05 0 2.7251e-05 5 2.75e-05 5   2.7501e-05 0 2.775e-05 0 2.7751e-05 5 2.8e-05 5   2.8001e-05 0 2.825e-05 0 2.8251e-05 5 2.85e-05 5   2.8501e-05 0 2.875e-05 0 2.8751e-05 5 2.9e-05 5   2.9001e-05 0 2.925e-05 0 2.9251e-05 5 2.95e-05 5   2.9501e-05 0 2.975e-05 0 2.9751e-05 5 3e-05 5   3.0001e-05 0 3.025e-05 0 3.0251e-05 5 3.05e-05 5   3.0501e-05 0 3.075e-05 0 3.0751e-05 5 3.1e-05 5   3.1001e-05 0 3.125e-05 0 3.1251e-05 5 3.15e-05 5   3.1501e-05 0 3.175e-05 0 3.1751e-05 5 3.2e-05 5   3.2001e-05 0 3.225e-05 0 3.2251e-05 5 3.25e-05 5   3.2501e-05 0 3.275e-05 0 3.2751e-05 5 3.3e-05 5   3.3001e-05 0 3.325e-05 0 3.3251e-05 5 3.35e-05 5   3.3501e-05 0 3.375e-05 0 3.3751e-05 5 3.4e-05 5   3.4001e-05 0 3.425e-05 0 3.4251e-05 5 3.45e-05 5   3.4501e-05 0 3.475e-05 0 3.4751e-05 5 3.5e-05 5   3.5001e-05 0 3.525e-05 0 3.5251e-05 5 3.55e-05 5   3.5501e-05 0 3.575e-05 0 3.5751e-05 5 3.6e-05 5   3.6001e-05 0 3.625e-05 0 3.6251e-05 5 3.65e-05 5   3.6501e-05 0 3.675e-05 0 3.6751e-05 5 3.7e-05 5   3.7001e-05 0 3.725e-05 0 3.7251e-05 5 3.75e-05 5   3.7501e-05 0 3.775e-05 0 3.7751e-05 5 3.8e-05 5   3.8001e-05 0 3.825e-05 0 3.8251e-05 5 3.85e-05 5   3.8501e-05 0 3.875e-05 0 3.8751e-05 5 3.9e-05 5   3.9001e-05 0 3.925e-05 0 3.9251e-05 5 3.95e-05 5   3.9501e-05 0 3.975e-05 0 3.9751e-05 5 4e-05 5   4.0001e-05 0 4.025e-05 0 )
V441 441 0 pwl (0 0 5e-07 0 5.01e-07 5 1e-06 5   1.001e-06 0 1.5e-06 0 1.501e-06 5 2e-06 5   2.001e-06 0 2.5e-06 0 2.501e-06 5 3e-06 5   3.001e-06 0 3.5e-06 0 3.501e-06 5 4e-06 5   4.001e-06 0 4.5e-06 0 4.501e-06 5 5e-06 5   5.001e-06 0 5.5e-06 0 5.501e-06 5 6e-06 5   6.001e-06 0 6.5e-06 0 6.501e-06 5 7e-06 5   7.001e-06 0 7.5e-06 0 7.501e-06 5 8e-06 5   8.001e-06 0 8.5e-06 0 8.501e-06 5 9e-06 5   9.001e-06 0 9.5e-06 0 9.501e-06 5 1e-05 5   1.0001e-05 0 1.05e-05 0 1.0501e-05 5 1.1e-05 5   1.1001e-05 0 1.15e-05 0 1.1501e-05 5 1.2e-05 5   1.2001e-05 0 1.25e-05 0 1.2501e-05 5 1.3e-05 5   1.3001e-05 0 1.35e-05 0 1.3501e-05 5 1.4e-05 5   1.4001e-05 0 1.45e-05 0 1.4501e-05 5 1.5e-05 5   1.5001e-05 0 1.55e-05 0 1.5501e-05 5 1.6e-05 5   1.6001e-05 0 1.65e-05 0 1.6501e-05 5 1.7e-05 5   1.7001e-05 0 1.75e-05 0 1.7501e-05 5 1.8e-05 5   1.8001e-05 0 1.85e-05 0 1.8501e-05 5 1.9e-05 5   1.9001e-05 0 1.95e-05 0 1.9501e-05 5 2e-05 5   2.0001e-05 0 2.05e-05 0 2.0501e-05 5 2.1e-05 5   2.1001e-05 0 2.15e-05 0 2.1501e-05 5 2.2e-05 5   2.2001e-05 0 2.25e-05 0 2.2501e-05 5 2.3e-05 5   2.3001e-05 0 2.35e-05 0 2.3501e-05 5 2.4e-05 5   2.4001e-05 0 2.45e-05 0 2.4501e-05 5 2.5e-05 5   2.5001e-05 0 2.55e-05 0 2.5501e-05 5 2.6e-05 5   2.6001e-05 0 2.65e-05 0 2.6501e-05 5 2.7e-05 5   2.7001e-05 0 2.75e-05 0 2.7501e-05 5 2.8e-05 5   2.8001e-05 0 2.85e-05 0 2.8501e-05 5 2.9e-05 5   2.9001e-05 0 2.95e-05 0 2.9501e-05 5 3e-05 5   3.0001e-05 0 3.05e-05 0 3.0501e-05 5 3.1e-05 5   3.1001e-05 0 3.15e-05 0 3.1501e-05 5 3.2e-05 5   3.2001e-05 0 3.25e-05 0 3.2501e-05 5 3.3e-05 5   3.3001e-05 0 3.35e-05 0 3.3501e-05 5 3.4e-05 5   3.4001e-05 0 3.45e-05 0 3.4501e-05 5 3.5e-05 5   3.5001e-05 0 3.55e-05 0 3.5501e-05 5 3.6e-05 5   3.6001e-05 0 3.65e-05 0 3.6501e-05 5 3.7e-05 5   3.7001e-05 0 3.75e-05 0 3.7501e-05 5 3.8e-05 5   3.8001e-05 0 3.85e-05 0 3.8501e-05 5 3.9e-05 5   3.9001e-05 0 3.95e-05 0 3.9501e-05 5 4e-05 5   4.0001e-05 0 4.05e-05 0 )
V442 442 0 pwl (0 0 1e-06 0 1.001e-06 5 2e-06 5   2.001e-06 0 3e-06 0 3.001e-06 5 4e-06 5   4.001e-06 0 5e-06 0 5.001e-06 5 6e-06 5   6.001e-06 0 7e-06 0 7.001e-06 5 8e-06 5   8.001e-06 0 9e-06 0 9.001e-06 5 1e-05 5   1.0001e-05 0 1.1e-05 0 1.1001e-05 5 1.2e-05 5   1.2001e-05 0 1.3e-05 0 1.3001e-05 5 1.4e-05 5   1.4001e-05 0 1.5e-05 0 1.5001e-05 5 1.6e-05 5   1.6001e-05 0 1.7e-05 0 1.7001e-05 5 1.8e-05 5   1.8001e-05 0 1.9e-05 0 1.9001e-05 5 2e-05 5   2.0001e-05 0 2.1e-05 0 2.1001e-05 5 2.2e-05 5   2.2001e-05 0 2.3e-05 0 2.3001e-05 5 2.4e-05 5   2.4001e-05 0 2.5e-05 0 2.5001e-05 5 2.6e-05 5   2.6001e-05 0 2.7e-05 0 2.7001e-05 5 2.8e-05 5   2.8001e-05 0 2.9e-05 0 2.9001e-05 5 3e-05 5   3.0001e-05 0 3.1e-05 0 3.1001e-05 5 3.2e-05 5   3.2001e-05 0 3.3e-05 0 3.3001e-05 5 3.4e-05 5   3.4001e-05 0 3.5e-05 0 3.5001e-05 5 3.6e-05 5   3.6001e-05 0 3.7e-05 0 3.7001e-05 5 3.8e-05 5   3.8001e-05 0 3.9e-05 0 3.9001e-05 5 4e-05 5   4.0001e-05 0 )
.print TRAN v(220) v(221) v(222) v(223) v(224) v(440) v(445) v(444) 
.options acct
.TRAN 1e-07 3e-05
.end
