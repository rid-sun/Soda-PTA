MOSAMP1 - MOS AMPLIFIER - DC/AC
*.OPTIONS ACCT  ABSTOL=10N VNTOL=10N
*.DC VIN -60MV +6MV 0.66MV
*.OP
*.AC DEC 10 100 10MEG
M1  15 15  1 32 M W=88.9U  L=25.4U
M2   1  1  2 32 M W=12.7U  L=266.7U
M3   2  2 30 32 M W=88.9U  L=25.4U
M4  15  5  4 32 M W=12.7U  L=106.7U
M5   4  4 30 32 M W=88.9U  L=12.7U
M6  15 15  5 32 M W=44.5U  L=25.4U
M7   5  0  8 32 M W=482.6U L=12.7U
M8   8  2 30 32 M W=88.9U  L=25.4U
M9  15 15  6 32 M W=44.5U  L=25.4U
M10  6 21  8 32 M W=482.6U L=12.7U
M11 15  6  7 32 M W=12.7U  L=106.7U
M12  7  4 30 32 M W=88.9U  L=12.7U
M13 15 10  9 32 M W=139.7U L=12.7U
M14  9 11 30 32 M W=139.7U L=12.7U
M15 15 15 12 32 M W=12.7U  L=207.8U
M16 12 12 11 32 M W=54.1U  L=12.7U
M17 11 11 30 32 M W=54.1U  L=12.7U
M18 15 15 10 32 M W=12.7U  L=45.2U
M19 10 12 13 32 M W=270.5U L=12.7U
M20 13  7 30 32 M W=270.5U L=12.7U
M21 15 10 14 32 M W=254U   L=12.7U
M22 14 11 30 32 M W=241.3U L=12.7U
M23 15 20 16 32 M W=19U    L=38.1U
M24 16 14 30 32 M W=406.4U L=12.7U
M25 15 15 20 32 M W=38.1U  L=42.7U
M26 20 16 30 32 M W=381U   L=25.4U
M27 20 15 66 32 M W=22.9U  L=7.6U
CC 7 9 40PF
CL 66 0 70PF
VIN 21 0 DC -30MV AC 1
VCCP 15 0 DC +15
VCCN 30 0 DC -15
VB 32 0 DC -20
.MODEL M NMOS(NSUB=2.2E15 UO=575 UCRIT=49K UEXP=0.1 TOX=0.11U XJ=2.95U    LEVEL=2 CGSO=1.5N CGDO=1.5N CBD=4.5F CBS=4.5F LD=2.4485U NSS=3.2E10)
*.PLOT DC V(20)
*.PRINT AC VDB(20) VP(20) VDB(66) VP(66)
*.PLOT  AC VDB(20) VP(20) VDB(66) VP(66)
*.END

.OPTIONS DELMAX=1000ns
.op
*.pstran convval=1.0e-05 initstep=1.0e-05 minstep=1.0e-06 maxstep=1.0e6 tau=1.0e-04 vbe0=0.0 kvgs0=0.0  tauramp=0.0
.end  