pchip.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.62249   kp = 6.32664e-05   gamma = 0.639243
+   phi = 0.31
+
+   cgso = 2.89e-10   cgdo = 2.89e-10
+   rsh = 60   cj = 0.000327
+   mj = 1.067   cjsw = 1.74e-10   mjsw = 0.195
+   tox = 2.25e-08   nsub = 1.066e+16
+   nss = 3e+10   nfs = 4.55168e+12   tpg = 1
+   xj = 9e-07   ld = 0   uo = 1215.74
+   ucrit = 174667   uexp = 0.0461235
+   vmax = 177269   neff = 4.6883
+
+   delta = 0
.model penh pmos
+ level = 2
+   vto = -0.63025   kp = 2.63544e-05   gamma = 0.618101
+   phi = 0.541111
+
+   cgso = 3.35e-10   cgdo = 3.35e-10
+   rsh = 150   cj = 0.000475
+   mj = 0.341   cjsw = 2.23e-10   mjsw = 0.307
+   tox = 2.25e-08   nsub = 6.57544e+16
+   nss = 3e+10   nfs = 1.66844e+11   tpg = -1
+   xj = 1.12799e-07   ld = 3e-08   uo = 361.941
+   ucrit = 637449   uexp = 0.0888696
+   vmax = 63253.3   neff = 0.64354
+
+   delta = 0
.subckt i 1 2 3 4 5
md1 2 7 6 2 nenh l=3e-06 w=4.5e-05 
+ as=3.375e-10 ad=2.41014e-09 ps=6e-05 pd=0.000160714 
+ nrs=0.166667 nrd=1.1902 
md2 3 7 6 3 penh l=3e-06 w=6.3e-05 
+ as=4.725e-10 ad=4.725e-10 ps=7.8e-05 pd=7.26921e-05 
+ nrs=0.119048 nrd=0.119048 
md3 7 5 2 2 nenh l=6e-06 w=4.5e-05 
+ as=2.41014e-09 ad=3.375e-10 ps=0.000160714 pd=6e-05 
+ nrs=1.1902 nrd=0.166667 
md4 7 5 3 3 penh l=6e-06 w=6.3e-05 
+ as=4.725e-10 ad=4.725e-10 ps=7.26921e-05 pd=7.8e-05 
+ nrs=0.119048 nrd=0.119048 
md5 2 2 5 2 nenh l=6e-06 w=6e-05 
+ as=2.5992e-08 ad=3.21353e-09 ps=0.001164 pd=0.000214285 
+ nrs=7.21999 nrd=0.892646 
md6 8 6 2 2 nenh l=3e-06 w=0.0001035 
+ as=5.54333e-09 ad=7.7625e-10 ps=0.000369643 pd=0.0001185 
+ nrs=0.517475 nrd=0.0724638 
md7 8 6 3 3 penh l=3e-06 w=0.000132 
+ as=9.9e-10 ad=9.9e-10 ps=0.000152308 pd=0.000147 
+ nrs=0.0568181 nrd=0.0568181 
md8 2 8 4 2 nenh l=3e-06 w=0.0001035 
+ as=7.7625e-10 ad=5.54333e-09 ps=0.0001185 pd=0.000369643 
+ nrs=0.0724638 nrd=0.517475 
md9 3 8 4 3 penh l=3e-06 w=0.000132 
+ as=9.9e-10 ad=9.9e-10 ps=0.000147 pd=0.000152308 
+ nrs=0.0568181 nrd=0.0568181 
c1 2 4 3.66898e-17
c2 2 8 3.86898e-17
c3 2 5 2.1064e-15
c4 2 7 1.47999e-17
c5 2 6 2.17999e-17
.ends i
.subckt four 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28
md10 29 30 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.44e-10 ps=2.75217e-05 pd=5.4e-05 
+ nrs=2.58877 nrd=4 
md11 31 32 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.44e-10 ps=2.75217e-05 pd=5.4e-05 
+ nrs=2.58877 nrd=4 
md12 28 34 33 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md13 28 36 35 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md14 28 38 37 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md15 39 40 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.215e-10 ps=2.75217e-05 pd=4.65e-05 
+ nrs=2.58877 nrd=3.375 
md16 41 42 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.215e-10 ps=2.75217e-05 pd=4.65e-05 
+ nrs=2.58877 nrd=3.375 
md17 28 44 43 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md18 28 46 45 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md19 28 48 47 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md20 49 50 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md21 51 52 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md22 24 53 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md23 23 54 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md24 28 56 55 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md25 57 58 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.2375e-10 ps=2.75217e-05 pd=4.725e-05 
+ nrs=2.58877 nrd=3.4375 
md26 59 60 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.2375e-10 ps=2.75217e-05 pd=4.725e-05 
+ nrs=2.58877 nrd=3.4375 
md27 28 62 61 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md28 28 64 63 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.71875 nrd=2.58877 
md29 28 11 65 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.71875 nrd=2.58877 
md30 66 67 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.484e-10 ps=5.50434e-05 pd=6.24e-05 
+ nrs=1.29438 nrd=1.725 
md31 28 69 68 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=9.31956e-11 ps=2.55e-05 pd=2.75217e-05 
+ nrs=2.09375 nrd=2.58877 
md32 70 71 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.484e-10 ps=5.50434e-05 pd=6.24e-05 
+ nrs=1.29438 nrd=1.725 
md33 28 6 72 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=9.31956e-11 ps=2.55e-05 pd=2.75217e-05 
+ nrs=2.09375 nrd=2.58877 
md34 73 74 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md35 75 76 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md36 28 78 77 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md37 79 80 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.62286e-10 ps=5.50434e-05 pd=6.25714e-05 
+ nrs=1.29438 nrd=1.82143 
md38 28 21 81 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md39 22 20 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.62286e-10 ps=5.50434e-05 pd=6.25714e-05 
+ nrs=1.29438 nrd=1.82143 
md40 82 83 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md41 28 85 84 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md42 86 87 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md43 28 89 88 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md44 28 91 90 28 penh l=3e-06 w=6e-06 
+ as=1.35e-10 ad=9.31956e-11 ps=4.5e-05 pd=2.75217e-05 
+ nrs=3.75 nrd=2.58877 
md45 92 93 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.08e-10 ps=2.75217e-05 pd=4.2e-05 
+ nrs=2.58877 nrd=3 
md46 94 95 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.08e-10 ps=2.75217e-05 pd=4.2e-05 
+ nrs=2.58877 nrd=3 
md47 28 97 96 28 penh l=3e-06 w=6e-06 
+ as=1.35e-10 ad=9.31956e-11 ps=4.5e-05 pd=2.75217e-05 
+ nrs=3.75 nrd=2.58877 
md48 83 98 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md49 28 99 85 28 penh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=1.86391e-10 ps=3.6e-05 pd=5.50434e-05 
+ nrs=0.9375 nrd=1.29438 
md50 87 100 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md51 28 101 89 28 penh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=1.86391e-10 ps=3.6e-05 pd=5.50434e-05 
+ nrs=0.9375 nrd=1.29438 
md52 28 103 102 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=9.31956e-11 ps=3.45e-05 pd=2.75217e-05 
+ nrs=3.4375 nrd=2.58877 
md53 104 25 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=8.1e-11 ps=2.75217e-05 pd=3.3e-05 
+ nrs=2.58877 nrd=2.25 
md54 28 19 17 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=9.31956e-11 ps=3.45e-05 pd=2.75217e-05 
+ nrs=3.4375 nrd=2.58877 
md55 105 26 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=8.1e-11 ps=2.75217e-05 pd=3.3e-05 
+ nrs=2.58877 nrd=2.25 
md56 28 107 106 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md57 28 109 108 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md58 103 15 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.295e-10 ps=5.50434e-05 pd=6e-05 
+ nrs=1.29438 nrd=1.59375 
md59 16 110 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.295e-10 ps=5.50434e-05 pd=6e-05 
+ nrs=1.29438 nrd=1.59375 
md60 28 112 111 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md61 28 114 113 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md62 14 115 28 28 penh l=6e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.89e-10 ps=5.50434e-05 pd=4.5e-05 
+ nrs=1.29438 nrd=1.3125 
md63 13 116 28 28 penh l=6e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.89e-10 ps=5.50434e-05 pd=4.5e-05 
+ nrs=1.29438 nrd=1.3125 
md64 117 118 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md65 119 120 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md66 28 122 121 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md67 28 124 123 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md68 28 126 125 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md69 28 128 127 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md70 129 130 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md71 131 132 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md72 28 134 133 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md73 28 136 135 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md74 122 137 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.44e-10 ps=2.75217e-05 pd=5.4e-05 
+ nrs=2.58877 nrd=4 
md75 124 138 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.44e-10 ps=2.75217e-05 pd=5.4e-05 
+ nrs=2.58877 nrd=4 
md76 28 140 139 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md77 28 142 141 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md78 28 144 143 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md79 145 146 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.215e-10 ps=2.75217e-05 pd=4.65e-05 
+ nrs=2.58877 nrd=3.375 
md80 147 148 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.215e-10 ps=2.75217e-05 pd=4.65e-05 
+ nrs=2.58877 nrd=3.375 
md81 28 150 149 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md82 28 64 151 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md83 152 153 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md84 28 11 12 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md85 154 155 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md86 28 157 156 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md87 28 159 158 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md88 160 161 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md89 162 163 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md90 164 165 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md91 166 167 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.67428e-10 ps=5.50434e-05 pd=6.34285e-05 
+ nrs=1.29438 nrd=1.85714 
md92 28 169 168 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md93 170 171 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.2375e-10 ps=2.75217e-05 pd=4.725e-05 
+ nrs=2.58877 nrd=3.4375 
md94 172 173 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.2375e-10 ps=2.75217e-05 pd=4.725e-05 
+ nrs=2.58877 nrd=3.4375 
md95 28 175 174 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md96 28 177 176 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.71875 nrd=2.58877 
md97 28 179 178 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.71875 nrd=2.58877 
md98 180 181 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.484e-10 ps=5.50434e-05 pd=6.24e-05 
+ nrs=1.29438 nrd=1.725 
md99 28 183 182 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=9.31956e-11 ps=2.55e-05 pd=2.75217e-05 
+ nrs=2.09375 nrd=2.58877 
md100 184 185 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.484e-10 ps=5.50434e-05 pd=6.24e-05 
+ nrs=1.29438 nrd=1.725 
md101 28 187 186 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=9.31956e-11 ps=2.55e-05 pd=2.75217e-05 
+ nrs=2.09375 nrd=2.58877 
md102 188 189 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md103 190 191 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md104 28 193 192 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md105 194 195 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.62286e-10 ps=5.50434e-05 pd=6.25714e-05 
+ nrs=1.29438 nrd=1.82143 
md106 28 197 196 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md107 198 199 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.62286e-10 ps=5.50434e-05 pd=6.25714e-05 
+ nrs=1.29438 nrd=1.82143 
md108 200 201 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md109 28 203 202 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md110 204 205 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md111 28 207 206 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md112 28 209 208 28 penh l=3e-06 w=6e-06 
+ as=1.35e-10 ad=9.31956e-11 ps=4.5e-05 pd=2.75217e-05 
+ nrs=3.75 nrd=2.58877 
md113 210 211 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.08e-10 ps=2.75217e-05 pd=4.2e-05 
+ nrs=2.58877 nrd=3 
md114 212 213 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=1.08e-10 ps=2.75217e-05 pd=4.2e-05 
+ nrs=2.58877 nrd=3 
md115 28 215 214 28 penh l=3e-06 w=6e-06 
+ as=1.35e-10 ad=9.31956e-11 ps=4.5e-05 pd=2.75217e-05 
+ nrs=3.75 nrd=2.58877 
md116 28 69 64 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md117 216 69 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md118 153 69 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md119 28 6 11 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md120 10 6 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md121 155 6 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md122 201 217 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md123 28 218 203 28 penh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=1.86391e-10 ps=3.6e-05 pd=5.50434e-05 
+ nrs=0.9375 nrd=1.29438 
md124 205 219 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.71e-10 ps=5.50434e-05 pd=4.2e-05 
+ nrs=1.29438 nrd=1.1875 
md125 28 220 207 28 penh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=1.86391e-10 ps=3.6e-05 pd=5.50434e-05 
+ nrs=0.9375 nrd=1.29438 
md126 221 222 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.1875e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.71875 
md127 223 222 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.0875e-11 ps=2.75217e-05 pd=2.4e-05 
+ nrs=2.58877 nrd=1.96875 
md128 224 4 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.1875e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.71875 
md129 225 4 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.0875e-11 ps=2.75217e-05 pd=2.4e-05 
+ nrs=2.58877 nrd=1.96875 
md130 28 227 226 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=9.31956e-11 ps=3.45e-05 pd=2.75217e-05 
+ nrs=3.4375 nrd=2.58877 
md131 228 229 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=8.1e-11 ps=2.75217e-05 pd=3.3e-05 
+ nrs=2.58877 nrd=2.25 
md132 28 9 230 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=9.31956e-11 ps=3.45e-05 pd=2.75217e-05 
+ nrs=3.4375 nrd=2.58877 
md133 231 232 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=8.1e-11 ps=2.75217e-05 pd=3.3e-05 
+ nrs=2.58877 nrd=2.25 
md134 28 233 118 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md135 28 234 120 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md136 227 235 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.295e-10 ps=5.50434e-05 pd=6e-05 
+ nrs=1.29438 nrd=1.59375 
md137 8 236 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=2.295e-10 ps=5.50434e-05 pd=6e-05 
+ nrs=1.29438 nrd=1.59375 
md138 28 177 130 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md139 237 238 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md140 28 179 132 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md141 239 240 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md142 28 183 177 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md143 241 183 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md144 238 183 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md145 28 187 179 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md146 242 187 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md147 240 187 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md148 243 244 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.1875e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.71875 
md149 245 244 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.0875e-11 ps=2.75217e-05 pd=2.4e-05 
+ nrs=2.58877 nrd=1.96875 
md150 246 247 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.1875e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.71875 
md151 248 247 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.0875e-11 ps=2.75217e-05 pd=2.4e-05 
+ nrs=2.58877 nrd=1.96875 
md152 28 250 249 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md153 28 252 251 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md154 28 254 253 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md155 28 1 183 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.31956e-11 ps=3e-05 pd=2.75217e-05 
+ nrs=2 nrd=2.58877 
md156 28 256 255 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md157 28 1 187 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.31956e-11 ps=3e-05 pd=2.75217e-05 
+ nrs=2 nrd=2.58877 
md158 28 257 254 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md159 244 2 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md160 252 257 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md161 28 258 256 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md162 247 2 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md163 250 258 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md164 28 260 259 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md165 28 262 261 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md166 28 264 263 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md167 28 1 69 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.31956e-11 ps=3e-05 pd=2.75217e-05 
+ nrs=2 nrd=2.58877 
md168 28 5 7 28 penh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=1.86391e-10 ps=4.2e-05 pd=5.50434e-05 
+ nrs=1.1875 nrd=1.29438 
md169 28 1 6 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.31956e-11 ps=3e-05 pd=2.75217e-05 
+ nrs=2 nrd=2.58877 
md170 28 265 264 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md171 222 2 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md172 262 265 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md173 28 3 5 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=1.86391e-10 ps=3.9e-05 pd=5.50434e-05 
+ nrs=1.0625 nrd=1.29438 
md174 4 2 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md175 260 3 28 28 penh l=3e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.35e-10 ps=5.50434e-05 pd=3.6e-05 
+ nrs=1.29438 nrd=0.9375 
md176 28 267 266 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md177 28 269 268 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md178 229 270 28 28 penh l=6e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.89e-10 ps=5.50434e-05 pd=4.5e-05 
+ nrs=1.29438 nrd=1.3125 
md179 232 271 28 28 penh l=6e-06 w=1.2e-05 
+ as=1.86391e-10 ad=1.89e-10 ps=5.50434e-05 pd=4.5e-05 
+ nrs=1.29438 nrd=1.3125 
md180 272 106 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md181 273 108 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=7.2e-11 ps=2.75217e-05 pd=3e-05 
+ nrs=2.58877 nrd=2 
md182 28 29 274 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md183 28 31 275 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.31956e-11 ps=2.1e-05 pd=2.75217e-05 
+ nrs=1.75 nrd=2.58877 
md184 28 277 276 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md185 28 279 278 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=1.86391e-10 ps=3.75e-05 pd=5.50434e-05 
+ nrs=1.5625 nrd=1.29438 
md186 280 151 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md187 281 12 28 28 penh l=3e-06 w=6e-06 
+ as=9.31956e-11 ad=6.3e-11 ps=2.75217e-05 pd=2.1e-05 
+ nrs=2.58877 nrd=1.75 
md188 28 283 282 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md189 28 285 284 28 penh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=9.31956e-11 ps=3.3e-05 pd=2.75217e-05 
+ nrs=2.75 nrd=2.58877 
md190 29 30 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.395e-10 ps=2.9923e-05 pd=6.09999e-05 
+ nrs=3.00641 nrd=3.875 
md191 31 32 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.395e-10 ps=2.9923e-05 pd=6.09999e-05 
+ nrs=3.00641 nrd=3.875 
md192 27 34 286 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md193 27 36 287 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md194 39 40 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.33875e-10 ps=2.9923e-05 pd=5.7e-05 
+ nrs=3.00641 nrd=3.71875 
md195 41 42 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.33875e-10 ps=2.9923e-05 pd=5.7e-05 
+ nrs=3.00641 nrd=3.71875 
md196 27 44 288 27 nenh l=3e-06 w=6e-06 
+ as=6.75e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=1.875 nrd=3.00641 
md197 27 38 289 27 nenh l=3e-06 w=6e-06 
+ as=6.75e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=1.875 nrd=3.00641 
md198 49 50 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md199 51 52 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md200 24 53 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md201 23 54 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md202 27 46 290 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md203 27 48 291 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md204 57 58 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.11375e-10 ps=2.9923e-05 pd=4.95e-05 
+ nrs=3.00641 nrd=3.09375 
md205 59 60 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.11375e-10 ps=2.9923e-05 pd=4.95e-05 
+ nrs=3.00641 nrd=3.09375 
md206 27 62 292 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md207 27 56 293 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md208 66 67 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.448e-10 ps=5.98461e-05 pd=7.55999e-05 
+ nrs=1.5032 nrd=1.7 
md209 70 71 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.448e-10 ps=5.98461e-05 pd=7.55999e-05 
+ nrs=1.5032 nrd=1.7 
md210 27 64 74 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md211 27 66 74 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md212 27 11 76 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md213 27 70 76 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md214 79 80 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.28857e-10 ps=5.98461e-05 pd=6.68571e-05 
+ nrs=1.5032 nrd=1.58928 
md215 22 20 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.28857e-10 ps=5.98461e-05 pd=6.68571e-05 
+ nrs=1.5032 nrd=1.58928 
md216 294 295 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md217 294 69 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md218 296 297 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md219 296 6 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md220 27 83 82 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md221 84 85 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md222 27 87 86 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md223 88 89 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md224 27 78 298 27 nenh l=3e-06 w=1.2e-05 
+ as=2.43e-10 ad=2.16461e-10 ps=5.4e-05 pd=5.98461e-05 
+ nrs=1.6875 nrd=1.5032 
md225 27 21 299 27 nenh l=3e-06 w=1.2e-05 
+ as=2.43e-10 ad=2.16461e-10 ps=5.4e-05 pd=5.98461e-05 
+ nrs=1.6875 nrd=1.5032 
md226 92 93 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.22625e-10 ps=2.9923e-05 pd=5.325e-05 
+ nrs=3.00641 nrd=3.40625 
md227 94 95 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.22625e-10 ps=2.9923e-05 pd=5.325e-05 
+ nrs=3.00641 nrd=3.40625 
md228 27 98 83 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md229 85 99 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md230 27 100 87 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md231 89 101 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md232 27 97 300 27 nenh l=3e-06 w=6e-06 
+ as=1.305e-10 ad=1.08231e-10 ps=4.95e-05 pd=2.9923e-05 
+ nrs=3.625 nrd=3.00641 
md233 27 91 301 27 nenh l=3e-06 w=6e-06 
+ as=1.305e-10 ad=1.08231e-10 ps=4.95e-05 pd=2.9923e-05 
+ nrs=3.625 nrd=3.00641 
md234 27 294 302 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md235 27 74 302 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md236 27 296 18 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md237 27 76 18 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md238 27 103 102 27 nenh l=3e-06 w=6e-06 
+ as=9.45e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=2.625 nrd=3.00641 
md239 104 25 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.485e-10 ps=5.98461e-05 pd=5.1e-05 
+ nrs=1.5032 nrd=1.03125 
md240 27 19 17 27 nenh l=3e-06 w=6e-06 
+ as=9.45e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=2.625 nrd=3.00641 
md241 105 26 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.485e-10 ps=5.98461e-05 pd=5.1e-05 
+ nrs=1.5032 nrd=1.03125 
md242 106 107 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md243 108 109 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md244 103 15 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.835e-10 ps=5.98461e-05 pd=7.8e-05 
+ nrs=1.5032 nrd=1.96875 
md245 16 110 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.835e-10 ps=5.98461e-05 pd=7.8e-05 
+ nrs=1.5032 nrd=1.96875 
md246 14 115 27 27 nenh l=6e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.89e-10 ps=5.98461e-05 pd=4.5e-05 
+ nrs=1.5032 nrd=1.3125 
md247 13 116 27 27 nenh l=6e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.89e-10 ps=5.98461e-05 pd=4.5e-05 
+ nrs=1.5032 nrd=1.3125 
md248 303 112 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md249 303 304 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md250 305 114 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md251 305 306 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md252 27 118 117 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md253 27 120 119 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md254 27 130 304 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md255 27 307 304 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md256 112 238 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md257 112 122 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md258 27 132 306 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md259 27 308 306 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md260 114 240 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md261 114 124 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md262 27 126 309 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md263 27 128 310 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md264 27 136 311 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md265 27 134 312 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md266 122 137 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.395e-10 ps=2.9923e-05 pd=6.09999e-05 
+ nrs=3.00641 nrd=3.875 
md267 124 138 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.395e-10 ps=2.9923e-05 pd=6.09999e-05 
+ nrs=3.00641 nrd=3.875 
md268 27 140 313 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md269 27 142 314 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md270 145 146 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.33875e-10 ps=2.9923e-05 pd=5.7e-05 
+ nrs=3.00641 nrd=3.71875 
md271 147 148 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.33875e-10 ps=2.9923e-05 pd=5.7e-05 
+ nrs=3.00641 nrd=3.71875 
md272 27 150 315 27 nenh l=3e-06 w=6e-06 
+ as=6.75e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=1.875 nrd=3.00641 
md273 27 144 316 27 nenh l=3e-06 w=6e-06 
+ as=6.75e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=1.875 nrd=3.00641 
md274 151 64 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md275 27 153 152 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md276 12 11 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md277 27 155 154 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md278 160 161 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md279 162 163 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md280 164 165 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md281 166 167 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.39143e-10 ps=5.98461e-05 pd=6.85713e-05 
+ nrs=1.5032 nrd=1.66071 
md282 27 157 317 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md283 27 159 318 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md284 170 171 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.11375e-10 ps=2.9923e-05 pd=4.95e-05 
+ nrs=3.00641 nrd=3.09375 
md285 172 173 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.11375e-10 ps=2.9923e-05 pd=4.95e-05 
+ nrs=3.00641 nrd=3.09375 
md286 27 175 319 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md287 27 169 320 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md288 180 181 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.448e-10 ps=5.98461e-05 pd=7.55999e-05 
+ nrs=1.5032 nrd=1.7 
md289 184 185 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.448e-10 ps=5.98461e-05 pd=7.55999e-05 
+ nrs=1.5032 nrd=1.7 
md290 27 177 189 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md291 27 180 189 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md292 27 179 191 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md293 27 184 191 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md294 194 195 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.28857e-10 ps=5.98461e-05 pd=6.68571e-05 
+ nrs=1.5032 nrd=1.58928 
md295 198 199 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.28857e-10 ps=5.98461e-05 pd=6.68571e-05 
+ nrs=1.5032 nrd=1.58928 
md296 321 322 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md297 321 183 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md298 323 324 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md299 323 187 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md300 27 201 200 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md301 202 203 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md302 27 205 204 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md303 206 207 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md304 107 69 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md305 107 222 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md306 109 6 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md307 109 4 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md308 27 193 325 27 nenh l=3e-06 w=1.2e-05 
+ as=2.43e-10 ad=2.16461e-10 ps=5.4e-05 pd=5.98461e-05 
+ nrs=1.6875 nrd=1.5032 
md309 27 197 326 27 nenh l=3e-06 w=1.2e-05 
+ as=2.43e-10 ad=2.16461e-10 ps=5.4e-05 pd=5.98461e-05 
+ nrs=1.6875 nrd=1.5032 
md310 210 211 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.22625e-10 ps=2.9923e-05 pd=5.325e-05 
+ nrs=3.00641 nrd=3.40625 
md311 212 213 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=1.22625e-10 ps=2.9923e-05 pd=5.325e-05 
+ nrs=3.00641 nrd=3.40625 
md312 64 69 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md313 27 69 216 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=1.08231e-10 ps=3.9e-05 pd=2.9923e-05 
+ nrs=2.75 nrd=3.00641 
md314 27 69 153 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md315 11 6 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md316 27 6 10 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=1.08231e-10 ps=3.9e-05 pd=2.9923e-05 
+ nrs=2.75 nrd=3.00641 
md317 27 6 155 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md318 27 217 201 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md319 203 218 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md320 27 219 205 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md321 207 220 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md322 27 215 327 27 nenh l=3e-06 w=6e-06 
+ as=1.305e-10 ad=1.08231e-10 ps=4.95e-05 pd=2.9923e-05 
+ nrs=3.625 nrd=3.00641 
md323 27 209 328 27 nenh l=3e-06 w=6e-06 
+ as=1.305e-10 ad=1.08231e-10 ps=4.95e-05 pd=2.9923e-05 
+ nrs=3.625 nrd=3.00641 
md324 27 321 329 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md325 27 189 329 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md326 27 323 330 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md327 27 191 330 27 nenh l=3e-06 w=6e-06 
+ as=9.59999e-11 ad=1.08231e-10 ps=3.79999e-05 pd=2.9923e-05 
+ nrs=2.66666 nrd=3.00641 
md328 27 227 226 27 nenh l=3e-06 w=6e-06 
+ as=9.45e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=2.625 nrd=3.00641 
md329 228 229 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.485e-10 ps=5.98461e-05 pd=5.1e-05 
+ nrs=1.5032 nrd=1.03125 
md330 27 9 230 27 nenh l=3e-06 w=6e-06 
+ as=9.45e-11 ad=1.08231e-10 ps=2.85e-05 pd=2.9923e-05 
+ nrs=2.625 nrd=3.00641 
md331 231 232 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.485e-10 ps=5.98461e-05 pd=5.1e-05 
+ nrs=1.5032 nrd=1.03125 
md332 118 233 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md333 120 234 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md334 227 235 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.835e-10 ps=5.98461e-05 pd=7.8e-05 
+ nrs=1.5032 nrd=1.96875 
md335 8 236 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.835e-10 ps=5.98461e-05 pd=7.8e-05 
+ nrs=1.5032 nrd=1.96875 
md336 130 177 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md337 27 238 237 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md338 132 179 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md339 27 240 239 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md340 233 183 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md341 233 244 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md342 234 187 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md343 234 247 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md344 177 183 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md345 27 183 241 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=1.08231e-10 ps=3.9e-05 pd=2.9923e-05 
+ nrs=2.75 nrd=3.00641 
md346 27 183 238 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md347 179 187 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.35e-10 ps=5.98461e-05 pd=3.6e-05 
+ nrs=1.5032 nrd=0.9375 
md348 27 187 242 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=1.08231e-10 ps=3.9e-05 pd=2.9923e-05 
+ nrs=2.75 nrd=3.00641 
md349 27 187 240 27 nenh l=3e-06 w=1.2e-05 
+ as=2.07e-10 ad=2.16461e-10 ps=4.8e-05 pd=5.98461e-05 
+ nrs=1.4375 nrd=1.5032 
md350 27 250 249 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md351 27 252 251 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md352 27 254 253 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md353 183 1 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md354 27 256 255 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md355 187 1 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md356 254 257 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.43e-10 ps=5.98461e-05 pd=5.4e-05 
+ nrs=1.5032 nrd=1.6875 
md357 27 2 244 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md358 27 257 252 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md359 256 258 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.43e-10 ps=5.98461e-05 pd=5.4e-05 
+ nrs=1.5032 nrd=1.6875 
md360 27 2 247 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md361 27 258 250 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md362 27 244 257 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md363 27 241 257 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md364 27 247 258 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md365 27 242 258 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md366 27 260 259 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md367 27 262 261 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md368 27 264 263 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md369 69 1 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md370 27 5 7 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md371 6 1 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md372 264 265 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.43e-10 ps=5.98461e-05 pd=5.4e-05 
+ nrs=1.5032 nrd=1.6875 
md373 27 2 222 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md374 27 265 262 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md375 5 3 27 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16461e-10 ad=2.43e-10 ps=5.98461e-05 pd=5.4e-05 
+ nrs=1.5032 nrd=1.6875 
md376 27 2 4 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md377 27 3 260 27 nenh l=3e-06 w=1.2e-05 
+ as=1.35e-10 ad=2.16461e-10 ps=3.6e-05 pd=5.98461e-05 
+ nrs=0.9375 nrd=1.5032 
md378 229 270 27 27 nenh l=6e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.89e-10 ps=5.98461e-05 pd=4.5e-05 
+ nrs=1.5032 nrd=1.3125 
md379 232 271 27 27 nenh l=6e-06 w=1.2e-05 
+ as=2.16461e-10 ad=1.89e-10 ps=5.98461e-05 pd=4.5e-05 
+ nrs=1.5032 nrd=1.3125 
md380 331 267 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md381 331 332 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md382 333 269 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md383 333 334 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=9e-11 ps=2.9923e-05 pd=3.6e-05 
+ nrs=3.00641 nrd=2.5 
md384 27 106 272 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md385 27 108 273 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md386 27 222 265 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md387 27 216 265 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md388 27 4 3 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md389 27 10 3 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md390 27 151 332 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md391 27 335 332 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md392 267 153 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md393 267 29 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md394 27 12 334 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md395 27 336 334 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md396 269 155 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md397 269 31 27 27 nenh l=3e-06 w=6e-06 
+ as=1.08231e-10 ad=7.2e-11 ps=2.9923e-05 pd=3e-05 
+ nrs=3.00641 nrd=2 
md398 27 277 337 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md399 27 279 338 27 nenh l=3e-06 w=1.2e-05 
+ as=1.71e-10 ad=2.16461e-10 ps=4.2e-05 pd=5.98461e-05 
+ nrs=1.1875 nrd=1.5032 
md400 27 285 339 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md401 27 283 340 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08231e-10 ps=3e-05 pd=2.9923e-05 
+ nrs=2 nrd=3.00641 
md402 341 83 29 27 nenh l=3e-06 w=6e-06 
+ as=1.395e-10 ad=8.69999e-11 ps=6.09999e-05 pd=3.1e-05 
+ nrs=3.875 nrd=2.41666 
md403 29 153 285 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.395e-10 ps=5.85e-05 pd=6.09999e-05 
+ nrs=4.375 nrd=3.875 
md404 29 82 341 28 penh l=3e-06 w=6e-06 
+ as=8.39999e-11 ad=1.44e-10 ps=3e-05 pd=5.4e-05 
+ nrs=2.33333 nrd=4 
md405 29 152 285 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.44e-10 ps=1.65e-05 pd=5.4e-05 
+ nrs=1.375 nrd=4 
md406 342 87 31 27 nenh l=3e-06 w=6e-06 
+ as=1.395e-10 ad=8.69999e-11 ps=6.09999e-05 pd=3.1e-05 
+ nrs=3.875 nrd=2.41666 
md407 31 155 283 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.395e-10 ps=5.85e-05 pd=6.09999e-05 
+ nrs=4.375 nrd=3.875 
md408 31 86 342 28 penh l=3e-06 w=6e-06 
+ as=8.39999e-11 ad=1.44e-10 ps=3e-05 pd=5.4e-05 
+ nrs=2.33333 nrd=4 
md409 31 154 283 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.44e-10 ps=1.65e-05 pd=5.4e-05 
+ nrs=1.375 nrd=4 
md410 339 262 30 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=7.2e-11 ps=4.2e-05 pd=3e-05 
+ nrs=3 nrd=2 
md411 284 261 30 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md412 340 260 32 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=7.2e-11 ps=4.2e-05 pd=3e-05 
+ nrs=3 nrd=2 
md413 282 259 32 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md414 33 263 50 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md415 35 7 53 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md416 286 264 50 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md417 49 64 34 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md418 34 263 51 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md419 49 151 34 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md420 34 264 51 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md421 335 85 341 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=7.65e-11 ps=3.1e-05 pd=2.55e-05 
+ nrs=2.41666 nrd=2.125 
md422 343 84 335 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.17e-10 ps=2.55e-05 pd=4.09999e-05 
+ nrs=2.125 nrd=3.25 
md423 341 84 335 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=8.39999e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.125 nrd=2.33333 
md424 335 85 343 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=7.65e-11 ps=4.2e-05 pd=2.55e-05 
+ nrs=3.33333 nrd=2.125 
md425 287 5 53 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md426 24 11 36 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md427 36 7 23 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md428 24 12 36 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md429 36 5 23 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md430 336 89 342 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=7.65e-11 ps=3.1e-05 pd=2.55e-05 
+ nrs=2.41666 nrd=2.125 
md431 344 88 336 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.17e-10 ps=2.55e-05 pd=4.09999e-05 
+ nrs=2.125 nrd=3.25 
md432 342 88 336 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=8.39999e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.125 nrd=2.33333 
md433 336 89 344 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=7.65e-11 ps=4.2e-05 pd=2.55e-05 
+ nrs=3.33333 nrd=2.125 
md434 37 259 42 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.9e-11 ps=3e-05 pd=3.3e-05 
+ nrs=2 nrd=2.75 
md435 39 82 341 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=1.33875e-10 ps=3.1e-05 pd=5.7e-05 
+ nrs=2.41666 nrd=3.71875 
md436 39 153 44 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.33875e-10 ps=5.85e-05 pd=5.7e-05 
+ nrs=4.375 nrd=3.71875 
md437 285 261 39 27 nenh l=3e-06 w=6e-06 
+ as=1.33875e-10 ad=1.575e-10 ps=5.7e-05 pd=5.85e-05 
+ nrs=3.71875 nrd=4.375 
md438 341 83 39 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=8.39999e-11 ps=4.65e-05 pd=3e-05 
+ nrs=3.375 nrd=2.33333 
md439 39 152 44 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.215e-10 ps=1.65e-05 pd=4.65e-05 
+ nrs=1.375 nrd=3.375 
md440 285 262 39 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=4.95e-11 ps=4.65e-05 pd=1.65e-05 
+ nrs=3.375 nrd=1.375 
md441 41 86 342 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=1.33875e-10 ps=3.1e-05 pd=5.7e-05 
+ nrs=2.41666 nrd=3.71875 
md442 41 155 38 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.33875e-10 ps=5.85e-05 pd=5.7e-05 
+ nrs=4.375 nrd=3.71875 
md443 283 259 41 27 nenh l=3e-06 w=6e-06 
+ as=1.33875e-10 ad=1.575e-10 ps=5.7e-05 pd=5.85e-05 
+ nrs=3.71875 nrd=4.375 
md444 342 87 41 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=8.39999e-11 ps=4.65e-05 pd=3e-05 
+ nrs=3.375 nrd=2.33333 
md445 41 154 38 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.215e-10 ps=1.65e-05 pd=4.65e-05 
+ nrs=1.375 nrd=3.375 
md446 283 260 41 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=4.95e-11 ps=4.65e-05 pd=1.65e-05 
+ nrs=3.375 nrd=1.375 
md447 43 261 40 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.9e-11 ps=3e-05 pd=3.3e-05 
+ nrs=2 nrd=2.75 
md448 343 83 57 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.17e-10 ps=4.95e-05 pd=4.09999e-05 
+ nrs=3.09375 nrd=3.25 
md449 92 82 343 27 nenh l=3e-06 w=6e-06 
+ as=1.17e-10 ad=1.22625e-10 ps=4.09999e-05 pd=5.325e-05 
+ nrs=3.25 nrd=3.40625 
md450 57 82 343 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=1.2375e-10 ps=4.2e-05 pd=4.725e-05 
+ nrs=3.33333 nrd=3.4375 
md451 343 83 92 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=1.2e-10 ps=4.2e-05 pd=4.2e-05 
+ nrs=3 nrd=3.33333 
md452 344 87 59 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.17e-10 ps=4.95e-05 pd=4.09999e-05 
+ nrs=3.09375 nrd=3.25 
md453 94 86 344 27 nenh l=3e-06 w=6e-06 
+ as=1.17e-10 ad=1.22625e-10 ps=4.09999e-05 pd=5.325e-05 
+ nrs=3.25 nrd=3.40625 
md454 59 86 344 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=1.2375e-10 ps=4.2e-05 pd=4.725e-05 
+ nrs=3.33333 nrd=3.4375 
md455 344 87 94 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=1.2e-10 ps=4.2e-05 pd=4.2e-05 
+ nrs=3 nrd=3.33333 
md456 44 261 57 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.575e-10 ps=4.95e-05 pd=5.85e-05 
+ nrs=3.09375 nrd=4.375 
md457 44 262 57 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=4.95e-11 ps=4.725e-05 pd=1.65e-05 
+ nrs=3.4375 nrd=1.375 
md458 288 262 40 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=6.75e-11 ps=4.2e-05 pd=2.85e-05 
+ nrs=3 nrd=1.875 
md459 38 259 59 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.575e-10 ps=4.95e-05 pd=5.85e-05 
+ nrs=3.09375 nrd=4.375 
md460 38 260 59 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=4.95e-11 ps=4.725e-05 pd=1.65e-05 
+ nrs=3.4375 nrd=1.375 
md461 289 260 42 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=6.75e-11 ps=4.2e-05 pd=2.85e-05 
+ nrs=3 nrd=1.875 
md462 45 263 52 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md463 49 82 345 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.19571e-10 ps=4.5e-05 pd=3.42856e-05 
+ nrs=3.58333 nrd=3.32143 
md464 295 85 345 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md465 345 83 66 27 nenh l=3e-06 w=6e-06 
+ as=1.224e-10 ad=1.29e-10 ps=3.77999e-05 pd=4.5e-05 
+ nrs=3.4 nrd=3.58333 
md466 345 83 49 28 penh l=3e-06 w=6e-06 
+ as=1.33714e-10 ad=1.26e-10 ps=3.17143e-05 pd=4.39999e-05 
+ nrs=3.71428 nrd=3.5 
md467 345 84 295 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md468 66 82 345 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.242e-10 ps=4.39999e-05 pd=3.12e-05 
+ nrs=3.5 nrd=3.45 
md469 346 83 51 27 nenh l=3e-06 w=6e-06 
+ as=1.19571e-10 ad=1.26e-10 ps=3.42856e-05 pd=4.39999e-05 
+ nrs=3.32143 nrd=3.5 
md470 346 84 295 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md471 79 82 346 27 nenh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.14428e-10 ps=4.39999e-05 pd=3.34285e-05 
+ nrs=3.5 nrd=3.17857 
md472 51 82 346 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.33714e-10 ps=4.5e-05 pd=3.17143e-05 
+ nrs=3.58333 nrd=3.71428 
md473 295 85 346 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md474 346 83 79 28 penh l=3e-06 w=6e-06 
+ as=1.31143e-10 ad=1.29e-10 ps=3.12857e-05 pd=4.5e-05 
+ nrs=3.64286 nrd=3.58333 
md475 47 7 54 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md476 24 86 347 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.19571e-10 ps=4.5e-05 pd=3.42856e-05 
+ nrs=3.58333 nrd=3.32143 
md477 297 89 347 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md478 347 87 70 27 nenh l=3e-06 w=6e-06 
+ as=1.224e-10 ad=1.29e-10 ps=3.77999e-05 pd=4.5e-05 
+ nrs=3.4 nrd=3.58333 
md479 347 87 24 28 penh l=3e-06 w=6e-06 
+ as=1.33714e-10 ad=1.26e-10 ps=3.17143e-05 pd=4.39999e-05 
+ nrs=3.71428 nrd=3.5 
md480 347 88 297 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md481 70 86 347 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.242e-10 ps=4.39999e-05 pd=3.12e-05 
+ nrs=3.5 nrd=3.45 
md482 348 87 23 27 nenh l=3e-06 w=6e-06 
+ as=1.19571e-10 ad=1.26e-10 ps=3.42856e-05 pd=4.39999e-05 
+ nrs=3.32143 nrd=3.5 
md483 348 88 297 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md484 22 86 348 27 nenh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.14428e-10 ps=4.39999e-05 pd=3.34285e-05 
+ nrs=3.5 nrd=3.17857 
md485 23 86 348 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.33714e-10 ps=4.5e-05 pd=3.17143e-05 
+ nrs=3.58333 nrd=3.71428 
md486 297 89 348 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md487 348 87 22 28 penh l=3e-06 w=6e-06 
+ as=1.31143e-10 ad=1.29e-10 ps=3.12857e-05 pd=4.5e-05 
+ nrs=3.64286 nrd=3.58333 
md488 277 263 49 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md489 277 264 49 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md490 51 64 46 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md491 51 151 46 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md492 279 7 24 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md493 279 5 24 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md494 23 11 48 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md495 23 12 48 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md496 290 264 52 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md497 46 263 79 27 nenh l=3e-06 w=1.2e-05 
+ as=2.28857e-10 ad=2.34e-10 ps=6.68571e-05 pd=5.25e-05 
+ nrs=1.58928 nrd=1.625 
md498 46 264 79 28 penh l=3e-06 w=1.2e-05 
+ as=2.62286e-10 ad=1.53e-10 ps=6.25714e-05 pd=2.55e-05 
+ nrs=1.82143 nrd=1.0625 
md499 291 5 54 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md500 48 7 22 27 nenh l=3e-06 w=1.2e-05 
+ as=2.28857e-10 ad=2.34e-10 ps=6.68571e-05 pd=5.25e-05 
+ nrs=1.58928 nrd=1.625 
md501 48 5 22 28 penh l=3e-06 w=1.2e-05 
+ as=2.62286e-10 ad=1.53e-10 ps=6.25714e-05 pd=2.55e-05 
+ nrs=1.82143 nrd=1.0625 
md502 55 259 60 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md503 57 153 62 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.11375e-10 ps=5.85e-05 pd=4.95e-05 
+ nrs=4.375 nrd=3.09375 
md504 57 152 62 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.2375e-10 ps=1.65e-05 pd=4.725e-05 
+ nrs=1.375 nrd=3.4375 
md505 59 155 56 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.11375e-10 ps=5.85e-05 pd=4.95e-05 
+ nrs=4.375 nrd=3.09375 
md506 59 154 56 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.2375e-10 ps=1.65e-05 pd=4.725e-05 
+ nrs=1.375 nrd=3.4375 
md507 61 261 58 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md508 62 261 92 27 nenh l=3e-06 w=6e-06 
+ as=1.22625e-10 ad=1.575e-10 ps=5.325e-05 pd=5.85e-05 
+ nrs=3.40625 nrd=4.375 
md509 62 262 92 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=4.95e-11 ps=4.2e-05 pd=1.65e-05 
+ nrs=3 nrd=1.375 
md510 292 262 58 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=7.2e-11 ps=3.9e-05 pd=3e-05 
+ nrs=2.75 nrd=2 
md511 56 259 94 27 nenh l=3e-06 w=6e-06 
+ as=1.22625e-10 ad=1.575e-10 ps=5.325e-05 pd=5.85e-05 
+ nrs=3.40625 nrd=4.375 
md512 56 260 94 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=4.95e-11 ps=4.2e-05 pd=1.65e-05 
+ nrs=3 nrd=1.375 
md513 293 260 60 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=7.2e-11 ps=3.9e-05 pd=3e-05 
+ nrs=2.75 nrd=2 
md514 74 66 63 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md515 76 70 65 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md516 66 64 277 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.448e-10 ps=5.25e-05 pd=7.55999e-05 
+ nrs=1.625 nrd=1.7 
md517 66 151 277 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.484e-10 ps=2.55e-05 pd=6.24e-05 
+ nrs=1.0625 nrd=1.725 
md518 294 295 68 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.09375 nrd=2 
md519 70 11 279 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.448e-10 ps=5.25e-05 pd=7.55999e-05 
+ nrs=1.625 nrd=1.7 
md520 70 12 279 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.484e-10 ps=2.55e-05 pd=6.24e-05 
+ nrs=1.0625 nrd=1.725 
md521 296 297 72 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.09375 nrd=2 
md522 302 294 73 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=8.1e-11 ps=2.1e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.25 
md523 18 296 75 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=8.1e-11 ps=2.1e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.25 
md524 77 263 80 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md525 79 64 78 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16e-10 ad=2.28857e-10 ps=4.95e-05 pd=6.68571e-05 
+ nrs=1.5 nrd=1.58928 
md526 79 151 78 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.62286e-10 ps=3.75e-05 pd=6.25714e-05 
+ nrs=1.5625 nrd=1.82143 
md527 81 7 20 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md528 22 11 21 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16e-10 ad=2.28857e-10 ps=4.95e-05 pd=6.68571e-05 
+ nrs=1.5 nrd=1.58928 
md529 22 12 21 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.62286e-10 ps=3.75e-05 pd=6.25714e-05 
+ nrs=1.5625 nrd=1.82143 
md530 298 264 80 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=2.43e-10 ps=6.6e-05 pd=5.4e-05 
+ nrs=2.1875 nrd=1.6875 
md531 78 263 102 27 nenh l=3e-06 w=1.2e-05 
+ as=1.89e-10 ad=2.16e-10 ps=5.7e-05 pd=4.95e-05 
+ nrs=1.3125 nrd=1.5 
md532 78 264 102 28 penh l=3e-06 w=1.2e-05 
+ as=2.475e-10 ad=2.25e-10 ps=6.9e-05 pd=3.75e-05 
+ nrs=1.71875 nrd=1.5625 
md533 299 5 20 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=2.43e-10 ps=6.6e-05 pd=5.4e-05 
+ nrs=2.1875 nrd=1.6875 
md534 21 7 17 27 nenh l=3e-06 w=1.2e-05 
+ as=1.89e-10 ad=2.16e-10 ps=5.7e-05 pd=4.95e-05 
+ nrs=1.3125 nrd=1.5 
md535 21 5 17 28 penh l=3e-06 w=1.2e-05 
+ as=2.475e-10 ad=2.25e-10 ps=6.9e-05 pd=3.75e-05 
+ nrs=1.71875 nrd=1.5625 
md536 90 259 95 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=1.35e-10 ps=2.7e-05 pd=4.5e-05 
+ nrs=1.75 nrd=3.75 
md537 92 153 97 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.22625e-10 ps=5.85e-05 pd=5.325e-05 
+ nrs=4.375 nrd=3.40625 
md538 92 152 97 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08e-10 ps=2.4e-05 pd=4.2e-05 
+ nrs=2 nrd=3 
md539 94 155 91 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.22625e-10 ps=5.85e-05 pd=5.325e-05 
+ nrs=4.375 nrd=3.40625 
md540 94 154 91 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08e-10 ps=2.4e-05 pd=4.2e-05 
+ nrs=2 nrd=3 
md541 96 261 93 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=1.35e-10 ps=2.7e-05 pd=4.5e-05 
+ nrs=1.75 nrd=3.75 
md542 97 261 104 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=1.575e-10 ps=2.55e-05 pd=5.85e-05 
+ nrs=2.0625 nrd=4.375 
md543 97 262 104 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=2.4e-05 
+ nrs=2.25 nrd=2 
md544 300 262 93 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.305e-10 ps=3e-05 pd=4.95e-05 
+ nrs=2 nrd=3.625 
md545 91 259 105 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=1.575e-10 ps=2.55e-05 pd=5.85e-05 
+ nrs=2.0625 nrd=4.375 
md546 91 260 105 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=2.4e-05 
+ nrs=2.25 nrd=2 
md547 301 260 95 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.305e-10 ps=3e-05 pd=4.95e-05 
+ nrs=2 nrd=3.625 
md548 102 107 98 27 nenh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=9.45e-11 ps=3.3e-05 pd=2.85e-05 
+ nrs=2.25 nrd=2.625 
md549 98 106 102 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=7.2e-11 ps=3.45e-05 pd=3e-05 
+ nrs=3.4375 nrd=2 
md550 99 107 104 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.0625 nrd=2 
md551 99 106 104 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md552 17 109 100 27 nenh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=9.45e-11 ps=3.3e-05 pd=2.85e-05 
+ nrs=2.25 nrd=2.625 
md553 100 108 17 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=7.2e-11 ps=3.45e-05 pd=3e-05 
+ nrs=3.4375 nrd=2 
md554 101 109 105 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.0625 nrd=2 
md555 101 108 105 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md556 302 106 110 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.59999e-11 ps=3e-05 pd=3.79999e-05 
+ nrs=2 nrd=2.66666 
md557 110 107 302 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md558 18 108 15 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.59999e-11 ps=3e-05 pd=3.79999e-05 
+ nrs=2 nrd=2.66666 
md559 15 109 18 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md560 111 304 303 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=6.3e-11 ps=4.8e-05 pd=2.1e-05 
+ nrs=3.5 nrd=1.75 
md561 113 306 305 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=6.3e-11 ps=4.8e-05 pd=2.1e-05 
+ nrs=3.5 nrd=1.75 
md562 116 120 305 27 nenh l=3e-06 w=6e-06 
+ as=9e-11 ad=8.1e-11 ps=3.6e-05 pd=3.3e-05 
+ nrs=2.5 nrd=2.25 
md563 116 119 305 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=8.1e-11 ps=4.8e-05 pd=3.3e-05 
+ nrs=3.5 nrd=2.25 
md564 115 118 303 27 nenh l=3e-06 w=6e-06 
+ as=9e-11 ad=8.1e-11 ps=3.6e-05 pd=3.3e-05 
+ nrs=2.5 nrd=2.25 
md565 115 117 303 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=8.1e-11 ps=4.8e-05 pd=3.3e-05 
+ nrs=3.5 nrd=2.25 
md566 121 238 112 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=6.3e-11 ps=3e-05 pd=2.1e-05 
+ nrs=2 nrd=1.75 
md567 123 240 114 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=6.3e-11 ps=3e-05 pd=2.1e-05 
+ nrs=2 nrd=1.75 
md568 125 253 181 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md569 127 255 185 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md570 304 307 129 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.75 nrd=2 
md571 306 308 131 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.75 nrd=2 
md572 309 254 181 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md573 126 253 160 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md574 180 177 126 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.448e-10 ps=5.25e-05 pd=7.55999e-05 
+ nrs=1.625 nrd=1.7 
md575 126 254 160 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md576 180 130 126 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.484e-10 ps=2.55e-05 pd=6.24e-05 
+ nrs=1.0625 nrd=1.725 
md577 310 256 185 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md578 128 255 164 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md579 184 179 128 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.448e-10 ps=5.25e-05 pd=7.55999e-05 
+ nrs=1.625 nrd=1.7 
md580 128 256 164 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md581 184 132 128 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.484e-10 ps=2.55e-05 pd=6.24e-05 
+ nrs=1.0625 nrd=1.725 
md582 133 249 138 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md583 135 251 137 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md584 122 238 136 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.395e-10 ps=5.85e-05 pd=6.09999e-05 
+ nrs=4.375 nrd=3.875 
md585 136 251 145 27 nenh l=3e-06 w=6e-06 
+ as=1.33875e-10 ad=1.575e-10 ps=5.7e-05 pd=5.85e-05 
+ nrs=3.71875 nrd=4.375 
md586 122 237 136 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.44e-10 ps=1.65e-05 pd=5.4e-05 
+ nrs=1.375 nrd=4 
md587 136 252 145 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=4.95e-11 ps=4.65e-05 pd=1.65e-05 
+ nrs=3.375 nrd=1.375 
md588 311 252 137 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=7.2e-11 ps=4.2e-05 pd=3e-05 
+ nrs=3 nrd=2 
md589 124 240 134 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.395e-10 ps=5.85e-05 pd=6.09999e-05 
+ nrs=4.375 nrd=3.875 
md590 134 249 147 27 nenh l=3e-06 w=6e-06 
+ as=1.33875e-10 ad=1.575e-10 ps=5.7e-05 pd=5.85e-05 
+ nrs=3.71875 nrd=4.375 
md591 124 239 134 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.44e-10 ps=1.65e-05 pd=5.4e-05 
+ nrs=1.375 nrd=4 
md592 134 250 147 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=4.95e-11 ps=4.65e-05 pd=1.65e-05 
+ nrs=3.375 nrd=1.375 
md593 312 250 138 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=7.2e-11 ps=4.2e-05 pd=3e-05 
+ nrs=3 nrd=2 
md594 349 201 122 27 nenh l=3e-06 w=6e-06 
+ as=1.395e-10 ad=8.69999e-11 ps=6.09999e-05 pd=3.1e-05 
+ nrs=3.875 nrd=2.41666 
md595 122 200 349 28 penh l=3e-06 w=6e-06 
+ as=8.39999e-11 ad=1.44e-10 ps=3e-05 pd=5.4e-05 
+ nrs=2.33333 nrd=4 
md596 350 205 124 27 nenh l=3e-06 w=6e-06 
+ as=1.395e-10 ad=8.69999e-11 ps=6.09999e-05 pd=3.1e-05 
+ nrs=3.875 nrd=2.41666 
md597 124 204 350 28 penh l=3e-06 w=6e-06 
+ as=8.39999e-11 ad=1.44e-10 ps=3e-05 pd=5.4e-05 
+ nrs=2.33333 nrd=4 
md598 139 253 161 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md599 141 255 165 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md600 313 254 161 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md601 160 177 140 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md602 140 253 162 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md603 160 130 140 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md604 140 254 162 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md605 307 203 349 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=7.65e-11 ps=3.1e-05 pd=2.55e-05 
+ nrs=2.41666 nrd=2.125 
md606 351 202 307 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.17e-10 ps=2.55e-05 pd=4.09999e-05 
+ nrs=2.125 nrd=3.25 
md607 349 202 307 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=8.39999e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.125 nrd=2.33333 
md608 307 203 351 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=7.65e-11 ps=4.2e-05 pd=2.55e-05 
+ nrs=3.33333 nrd=2.125 
md609 314 256 165 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md610 164 179 142 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md611 142 255 166 27 nenh l=3e-06 w=1.2e-05 
+ as=2.39143e-10 ad=2.34e-10 ps=6.85713e-05 pd=5.25e-05 
+ nrs=1.66071 nrd=1.625 
md612 164 132 142 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md613 142 256 166 28 penh l=3e-06 w=1.2e-05 
+ as=2.67428e-10 ad=1.53e-10 ps=6.34285e-05 pd=2.55e-05 
+ nrs=1.85714 nrd=1.0625 
md614 308 207 350 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=7.65e-11 ps=3.1e-05 pd=2.55e-05 
+ nrs=2.41666 nrd=2.125 
md615 352 206 308 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.17e-10 ps=2.55e-05 pd=4.09999e-05 
+ nrs=2.125 nrd=3.25 
md616 350 206 308 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=8.39999e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.125 nrd=2.33333 
md617 308 207 352 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=7.65e-11 ps=4.2e-05 pd=2.55e-05 
+ nrs=3.33333 nrd=2.125 
md618 143 249 148 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.9e-11 ps=3e-05 pd=3.3e-05 
+ nrs=2 nrd=2.75 
md619 145 200 349 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=1.33875e-10 ps=3.1e-05 pd=5.7e-05 
+ nrs=2.41666 nrd=3.71875 
md620 145 238 150 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.33875e-10 ps=5.85e-05 pd=5.7e-05 
+ nrs=4.375 nrd=3.71875 
md621 349 201 145 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=8.39999e-11 ps=4.65e-05 pd=3e-05 
+ nrs=3.375 nrd=2.33333 
md622 145 237 150 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.215e-10 ps=1.65e-05 pd=4.65e-05 
+ nrs=1.375 nrd=3.375 
md623 147 204 350 27 nenh l=3e-06 w=6e-06 
+ as=8.69999e-11 ad=1.33875e-10 ps=3.1e-05 pd=5.7e-05 
+ nrs=2.41666 nrd=3.71875 
md624 147 240 144 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.33875e-10 ps=5.85e-05 pd=5.7e-05 
+ nrs=4.375 nrd=3.71875 
md625 350 205 147 28 penh l=3e-06 w=6e-06 
+ as=1.215e-10 ad=8.39999e-11 ps=4.65e-05 pd=3e-05 
+ nrs=3.375 nrd=2.33333 
md626 147 239 144 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.215e-10 ps=1.65e-05 pd=4.65e-05 
+ nrs=1.375 nrd=3.375 
md627 149 251 146 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.9e-11 ps=3e-05 pd=3.3e-05 
+ nrs=2 nrd=2.75 
md628 351 201 170 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.17e-10 ps=4.95e-05 pd=4.09999e-05 
+ nrs=3.09375 nrd=3.25 
md629 210 200 351 27 nenh l=3e-06 w=6e-06 
+ as=1.17e-10 ad=1.22625e-10 ps=4.09999e-05 pd=5.325e-05 
+ nrs=3.25 nrd=3.40625 
md630 170 200 351 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=1.2375e-10 ps=4.2e-05 pd=4.725e-05 
+ nrs=3.33333 nrd=3.4375 
md631 351 201 210 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=1.2e-10 ps=4.2e-05 pd=4.2e-05 
+ nrs=3 nrd=3.33333 
md632 352 205 172 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.17e-10 ps=4.95e-05 pd=4.09999e-05 
+ nrs=3.09375 nrd=3.25 
md633 212 204 352 27 nenh l=3e-06 w=6e-06 
+ as=1.17e-10 ad=1.22625e-10 ps=4.09999e-05 pd=5.325e-05 
+ nrs=3.25 nrd=3.40625 
md634 172 204 352 28 penh l=3e-06 w=6e-06 
+ as=1.2e-10 ad=1.2375e-10 ps=4.2e-05 pd=4.725e-05 
+ nrs=3.33333 nrd=3.4375 
md635 352 205 212 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=1.2e-10 ps=4.2e-05 pd=4.2e-05 
+ nrs=3 nrd=3.33333 
md636 150 251 170 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.575e-10 ps=4.95e-05 pd=5.85e-05 
+ nrs=3.09375 nrd=4.375 
md637 150 252 170 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=4.95e-11 ps=4.725e-05 pd=1.65e-05 
+ nrs=3.4375 nrd=1.375 
md638 315 252 146 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=6.75e-11 ps=4.2e-05 pd=2.85e-05 
+ nrs=3 nrd=1.875 
md639 144 249 172 27 nenh l=3e-06 w=6e-06 
+ as=1.11375e-10 ad=1.575e-10 ps=4.95e-05 pd=5.85e-05 
+ nrs=3.09375 nrd=4.375 
md640 144 250 172 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=4.95e-11 ps=4.725e-05 pd=1.65e-05 
+ nrs=3.4375 nrd=1.375 
md641 316 250 148 27 nenh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=6.75e-11 ps=4.2e-05 pd=2.85e-05 
+ nrs=3 nrd=1.875 
md642 156 253 163 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md643 160 200 353 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.19571e-10 ps=4.5e-05 pd=3.42856e-05 
+ nrs=3.58333 nrd=3.32143 
md644 322 203 353 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md645 353 201 180 27 nenh l=3e-06 w=6e-06 
+ as=1.224e-10 ad=1.29e-10 ps=3.77999e-05 pd=4.5e-05 
+ nrs=3.4 nrd=3.58333 
md646 353 201 160 28 penh l=3e-06 w=6e-06 
+ as=1.33714e-10 ad=1.26e-10 ps=3.17143e-05 pd=4.39999e-05 
+ nrs=3.71428 nrd=3.5 
md647 353 202 322 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md648 180 200 353 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.242e-10 ps=4.39999e-05 pd=3.12e-05 
+ nrs=3.5 nrd=3.45 
md649 354 201 162 27 nenh l=3e-06 w=6e-06 
+ as=1.19571e-10 ad=1.26e-10 ps=3.42856e-05 pd=4.39999e-05 
+ nrs=3.32143 nrd=3.5 
md650 354 202 322 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md651 194 200 354 27 nenh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.14428e-10 ps=4.39999e-05 pd=3.34285e-05 
+ nrs=3.5 nrd=3.17857 
md652 162 200 354 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.33714e-10 ps=4.5e-05 pd=3.17143e-05 
+ nrs=3.58333 nrd=3.71428 
md653 322 203 354 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md654 354 201 194 28 penh l=3e-06 w=6e-06 
+ as=1.31143e-10 ad=1.29e-10 ps=3.12857e-05 pd=4.5e-05 
+ nrs=3.64286 nrd=3.58333 
md655 158 255 167 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md656 164 204 355 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.19571e-10 ps=4.5e-05 pd=3.42856e-05 
+ nrs=3.58333 nrd=3.32143 
md657 324 207 355 27 nenh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md658 355 205 184 27 nenh l=3e-06 w=6e-06 
+ as=1.224e-10 ad=1.29e-10 ps=3.77999e-05 pd=4.5e-05 
+ nrs=3.4 nrd=3.58333 
md659 355 205 164 28 penh l=3e-06 w=6e-06 
+ as=1.33714e-10 ad=1.26e-10 ps=3.17143e-05 pd=4.39999e-05 
+ nrs=3.71428 nrd=3.5 
md660 355 206 324 28 penh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md661 184 204 355 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.242e-10 ps=4.39999e-05 pd=3.12e-05 
+ nrs=3.5 nrd=3.45 
md662 356 205 166 27 nenh l=3e-06 w=6e-06 
+ as=1.19571e-10 ad=1.26e-10 ps=3.42856e-05 pd=4.39999e-05 
+ nrs=3.32143 nrd=3.5 
md663 356 206 324 27 nenh l=3e-06 w=6e-06 
+ as=7.65e-11 ad=1.26e-10 ps=2.55e-05 pd=4.39999e-05 
+ nrs=2.125 nrd=3.5 
md664 198 204 356 27 nenh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=1.14428e-10 ps=4.39999e-05 pd=3.34285e-05 
+ nrs=3.5 nrd=3.17857 
md665 166 204 356 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=1.33714e-10 ps=4.5e-05 pd=3.17143e-05 
+ nrs=3.58333 nrd=3.71428 
md666 324 207 356 28 penh l=3e-06 w=6e-06 
+ as=1.29e-10 ad=7.65e-11 ps=4.5e-05 pd=2.55e-05 
+ nrs=3.58333 nrd=2.125 
md667 356 205 198 28 penh l=3e-06 w=6e-06 
+ as=1.31143e-10 ad=1.29e-10 ps=3.12857e-05 pd=4.5e-05 
+ nrs=3.64286 nrd=3.58333 
md668 162 177 157 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md669 162 130 157 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md670 166 179 159 27 nenh l=3e-06 w=1.2e-05 
+ as=2.34e-10 ad=2.39143e-10 ps=5.25e-05 pd=6.85713e-05 
+ nrs=1.625 nrd=1.66071 
md671 166 132 159 28 penh l=3e-06 w=1.2e-05 
+ as=1.53e-10 ad=2.67428e-10 ps=2.55e-05 pd=6.34285e-05 
+ nrs=1.0625 nrd=1.85714 
md672 317 254 163 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md673 157 253 194 27 nenh l=3e-06 w=1.2e-05 
+ as=2.28857e-10 ad=2.34e-10 ps=6.68571e-05 pd=5.25e-05 
+ nrs=1.58928 nrd=1.625 
md674 157 254 194 28 penh l=3e-06 w=1.2e-05 
+ as=2.62286e-10 ad=1.53e-10 ps=6.25714e-05 pd=2.55e-05 
+ nrs=1.82143 nrd=1.0625 
md675 318 256 167 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md676 159 255 198 27 nenh l=3e-06 w=1.2e-05 
+ as=2.28857e-10 ad=2.34e-10 ps=6.68571e-05 pd=5.25e-05 
+ nrs=1.58928 nrd=1.625 
md677 159 256 198 28 penh l=3e-06 w=1.2e-05 
+ as=2.62286e-10 ad=1.53e-10 ps=6.25714e-05 pd=2.55e-05 
+ nrs=1.82143 nrd=1.0625 
md678 168 249 173 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md679 170 238 175 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.11375e-10 ps=5.85e-05 pd=4.95e-05 
+ nrs=4.375 nrd=3.09375 
md680 170 237 175 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.2375e-10 ps=1.65e-05 pd=4.725e-05 
+ nrs=1.375 nrd=3.4375 
md681 172 240 169 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.11375e-10 ps=5.85e-05 pd=4.95e-05 
+ nrs=4.375 nrd=3.09375 
md682 172 239 169 28 penh l=3e-06 w=6e-06 
+ as=4.95e-11 ad=1.2375e-10 ps=1.65e-05 pd=4.725e-05 
+ nrs=1.375 nrd=3.4375 
md683 174 251 171 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=9.9e-11 ps=2.7e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.75 
md684 175 251 210 27 nenh l=3e-06 w=6e-06 
+ as=1.22625e-10 ad=1.575e-10 ps=5.325e-05 pd=5.85e-05 
+ nrs=3.40625 nrd=4.375 
md685 175 252 210 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=4.95e-11 ps=4.2e-05 pd=1.65e-05 
+ nrs=3 nrd=1.375 
md686 319 252 171 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=7.2e-11 ps=3.9e-05 pd=3e-05 
+ nrs=2.75 nrd=2 
md687 169 249 212 27 nenh l=3e-06 w=6e-06 
+ as=1.22625e-10 ad=1.575e-10 ps=5.325e-05 pd=5.85e-05 
+ nrs=3.40625 nrd=4.375 
md688 169 250 212 28 penh l=3e-06 w=6e-06 
+ as=1.08e-10 ad=4.95e-11 ps=4.2e-05 pd=1.65e-05 
+ nrs=3 nrd=1.375 
md689 320 250 173 27 nenh l=3e-06 w=6e-06 
+ as=9.9e-11 ad=7.2e-11 ps=3.9e-05 pd=3e-05 
+ nrs=2.75 nrd=2 
md690 189 180 176 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md691 191 184 178 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md692 321 322 182 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.09375 nrd=2 
md693 323 324 186 28 penh l=3e-06 w=6e-06 
+ as=7.5375e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.09375 nrd=2 
md694 329 321 188 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=8.1e-11 ps=2.1e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.25 
md695 330 323 190 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=8.1e-11 ps=2.1e-05 pd=3.3e-05 
+ nrs=1.75 nrd=2.25 
md696 192 253 195 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md697 194 177 193 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16e-10 ad=2.28857e-10 ps=4.95e-05 pd=6.68571e-05 
+ nrs=1.5 nrd=1.58928 
md698 194 130 193 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.62286e-10 ps=3.75e-05 pd=6.25714e-05 
+ nrs=1.5625 nrd=1.82143 
md699 196 255 199 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md700 198 179 197 27 nenh l=3e-06 w=1.2e-05 
+ as=2.16e-10 ad=2.28857e-10 ps=4.95e-05 pd=6.68571e-05 
+ nrs=1.5 nrd=1.58928 
md701 198 132 197 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.62286e-10 ps=3.75e-05 pd=6.25714e-05 
+ nrs=1.5625 nrd=1.82143 
md702 223 69 107 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=7.0875e-11 ps=3e-05 pd=2.4e-05 
+ nrs=2 nrd=1.96875 
md703 225 6 109 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=7.0875e-11 ps=3e-05 pd=2.4e-05 
+ nrs=2 nrd=1.96875 
md704 325 254 195 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=2.43e-10 ps=6.6e-05 pd=5.4e-05 
+ nrs=2.1875 nrd=1.6875 
md705 193 253 226 27 nenh l=3e-06 w=1.2e-05 
+ as=1.89e-10 ad=2.16e-10 ps=5.7e-05 pd=4.95e-05 
+ nrs=1.3125 nrd=1.5 
md706 193 254 226 28 penh l=3e-06 w=1.2e-05 
+ as=2.475e-10 ad=2.25e-10 ps=6.9e-05 pd=3.75e-05 
+ nrs=1.71875 nrd=1.5625 
md707 326 256 199 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=2.43e-10 ps=6.6e-05 pd=5.4e-05 
+ nrs=2.1875 nrd=1.6875 
md708 197 255 230 27 nenh l=3e-06 w=1.2e-05 
+ as=1.89e-10 ad=2.16e-10 ps=5.7e-05 pd=4.95e-05 
+ nrs=1.3125 nrd=1.5 
md709 197 256 230 28 penh l=3e-06 w=1.2e-05 
+ as=2.475e-10 ad=2.25e-10 ps=6.9e-05 pd=3.75e-05 
+ nrs=1.71875 nrd=1.5625 
md710 208 249 213 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=1.35e-10 ps=2.7e-05 pd=4.5e-05 
+ nrs=1.75 nrd=3.75 
md711 210 238 215 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.22625e-10 ps=5.85e-05 pd=5.325e-05 
+ nrs=4.375 nrd=3.40625 
md712 210 237 215 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08e-10 ps=2.4e-05 pd=4.2e-05 
+ nrs=2 nrd=3 
md713 212 240 209 27 nenh l=3e-06 w=6e-06 
+ as=1.575e-10 ad=1.22625e-10 ps=5.85e-05 pd=5.325e-05 
+ nrs=4.375 nrd=3.40625 
md714 212 239 209 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.08e-10 ps=2.4e-05 pd=4.2e-05 
+ nrs=2 nrd=3 
md715 214 251 211 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=1.35e-10 ps=2.7e-05 pd=4.5e-05 
+ nrs=1.75 nrd=3.75 
md716 215 251 228 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=1.575e-10 ps=2.55e-05 pd=5.85e-05 
+ nrs=2.0625 nrd=4.375 
md717 215 252 228 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=2.4e-05 
+ nrs=2.25 nrd=2 
md718 327 252 211 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.305e-10 ps=3e-05 pd=4.95e-05 
+ nrs=2 nrd=3.625 
md719 209 249 231 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=1.575e-10 ps=2.55e-05 pd=5.85e-05 
+ nrs=2.0625 nrd=4.375 
md720 209 250 231 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=2.4e-05 
+ nrs=2.25 nrd=2 
md721 328 250 213 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=1.305e-10 ps=3e-05 pd=4.95e-05 
+ nrs=2 nrd=3.625 
md722 226 233 217 27 nenh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=9.45e-11 ps=3.3e-05 pd=2.85e-05 
+ nrs=2.25 nrd=2.625 
md723 217 118 226 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=7.2e-11 ps=3.45e-05 pd=3e-05 
+ nrs=3.4375 nrd=2 
md724 218 233 228 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.0625 nrd=2 
md725 218 118 228 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md726 230 234 219 27 nenh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=9.45e-11 ps=3.3e-05 pd=2.85e-05 
+ nrs=2.25 nrd=2.625 
md727 219 120 230 28 penh l=3e-06 w=6e-06 
+ as=1.2375e-10 ad=7.2e-11 ps=3.45e-05 pd=3e-05 
+ nrs=3.4375 nrd=2 
md728 220 234 231 27 nenh l=3e-06 w=6e-06 
+ as=7.425e-11 ad=7.2e-11 ps=2.55e-05 pd=3e-05 
+ nrs=2.0625 nrd=2 
md729 220 120 231 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md730 265 216 221 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md731 3 10 224 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md732 329 118 236 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.59999e-11 ps=3e-05 pd=3.79999e-05 
+ nrs=2 nrd=2.66666 
md733 236 233 329 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md734 330 120 235 27 nenh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=9.59999e-11 ps=3e-05 pd=3.79999e-05 
+ nrs=2 nrd=2.66666 
md735 235 234 330 28 penh l=3e-06 w=6e-06 
+ as=8.1e-11 ad=7.2e-11 ps=3.3e-05 pd=3e-05 
+ nrs=2.25 nrd=2 
md736 245 183 233 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=7.0875e-11 ps=3e-05 pd=2.4e-05 
+ nrs=2 nrd=1.96875 
md737 248 187 234 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=7.0875e-11 ps=3e-05 pd=2.4e-05 
+ nrs=2 nrd=1.96875 
md738 257 241 243 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md739 258 242 246 28 penh l=3e-06 w=6e-06 
+ as=6.1875e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.71875 nrd=2 
md740 266 332 331 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=6.3e-11 ps=4.8e-05 pd=2.1e-05 
+ nrs=3.5 nrd=1.75 
md741 268 334 333 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=6.3e-11 ps=4.8e-05 pd=2.1e-05 
+ nrs=3.5 nrd=1.75 
md742 271 108 333 27 nenh l=3e-06 w=6e-06 
+ as=9e-11 ad=8.1e-11 ps=3.6e-05 pd=3.3e-05 
+ nrs=2.5 nrd=2.25 
md743 271 273 333 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=8.1e-11 ps=4.8e-05 pd=3.3e-05 
+ nrs=3.5 nrd=2.25 
md744 270 106 331 27 nenh l=3e-06 w=6e-06 
+ as=9e-11 ad=8.1e-11 ps=3.6e-05 pd=3.3e-05 
+ nrs=2.5 nrd=2.25 
md745 270 272 331 28 penh l=3e-06 w=6e-06 
+ as=1.26e-10 ad=8.1e-11 ps=4.8e-05 pd=3.3e-05 
+ nrs=3.5 nrd=2.25 
md746 274 153 267 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=6.3e-11 ps=3e-05 pd=2.1e-05 
+ nrs=2 nrd=1.75 
md747 275 155 269 28 penh l=3e-06 w=6e-06 
+ as=7.2e-11 ad=6.3e-11 ps=3e-05 pd=2.1e-05 
+ nrs=2 nrd=1.75 
md748 276 263 67 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md749 278 7 71 28 penh l=3e-06 w=1.2e-05 
+ as=2.25e-10 ad=2.25e-10 ps=5.1e-05 pd=3.75e-05 
+ nrs=1.5625 nrd=1.5625 
md750 332 335 280 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.75 nrd=2 
md751 334 336 281 28 penh l=3e-06 w=6e-06 
+ as=6.3e-11 ad=7.2e-11 ps=2.1e-05 pd=3e-05 
+ nrs=1.75 nrd=2 
md752 337 264 67 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
md753 338 5 71 27 nenh l=3e-06 w=1.2e-05 
+ as=3.15e-10 ad=1.71e-10 ps=6.6e-05 pd=4.2e-05 
+ nrs=2.1875 nrd=1.1875 
c6 340 27 2.67999e-18
c7 283 27 1.51099e-17
c8 339 27 2.67999e-18
c9 285 27 1.51099e-17
c10 71 27 1.37899e-17
c11 67 27 1.37899e-17
c12 279 27 1.63299e-17
c13 338 27 3.19999e-18
c14 277 27 1.63299e-17
c15 337 27 3.19999e-18
c16 269 27 2.30199e-17
c17 334 27 2.40199e-17
c18 267 27 2.30199e-17
c19 332 27 2.40199e-17
c20 1 27 1.06199e-18
c21 3 27 6.50197e-17
c22 265 27 6.50197e-17
c23 273 27 1.11799e-17
c24 272 27 1.11799e-17
c25 333 27 1.51599e-17
c26 331 27 1.51599e-17
c27 270 27 5.29098e-17
c28 271 27 5.29098e-17
c29 232 27 7.63097e-17
c30 229 27 7.63097e-17
c31 260 27 1.28439e-16
c32 4 27 3.14399e-17
c33 5 27 1.29629e-16
c34 262 27 1.28439e-16
c35 222 27 3.14399e-17
c36 264 27 1.29629e-16
c37 6 27 1.23179e-16
c38 7 27 1.2202e-16
c39 69 27 1.23179e-16
c40 263 27 1.2202e-16
c41 261 27 1.1202e-16
c42 259 27 1.1202e-16
c43 258 27 6.50197e-17
c44 257 27 6.50197e-17
c45 250 27 1.28439e-16
c46 247 27 3.14399e-17
c47 256 27 1.29629e-16
c48 252 27 1.28439e-16
c49 244 27 3.14399e-17
c50 254 27 1.29629e-16
c51 187 27 1.23179e-16
c52 255 27 1.2202e-16
c53 183 27 1.23179e-16
c54 253 27 1.2202e-16
c55 251 27 1.1202e-16
c56 249 27 1.1202e-16
c57 240 27 1.42959e-16
c58 242 27 1.40799e-17
c59 179 27 1.44349e-16
c60 238 27 1.42959e-16
c61 241 27 1.40799e-17
c62 177 27 1.44349e-16
c63 234 27 6.30198e-17
c64 233 27 6.30198e-17
c65 239 27 8.39596e-17
c66 132 27 1.14349e-16
c67 237 27 8.39596e-17
c68 130 27 1.14349e-16
c69 236 27 5.11798e-17
c70 235 27 5.11798e-17
c71 8 27 2.59799e-17
c72 227 27 3.99799e-17
c73 120 27 1.39259e-16
c74 118 27 1.39259e-16
c75 231 27 3.44299e-17
c76 230 27 4.68198e-17
c77 228 27 3.44299e-17
c78 226 27 4.68198e-17
c79 330 27 2.74601e-17
c80 329 27 2.74601e-17
c81 213 27 1.37499e-17
c82 211 27 1.37499e-17
c83 220 27 2.11799e-17
c84 219 27 1.74799e-17
c85 218 27 2.11799e-17
c86 217 27 1.74799e-17
c87 328 27 2.57999e-18
c88 209 27 1.62599e-17
c89 327 27 2.57999e-18
c90 215 27 1.62599e-17
c91 207 27 8.24397e-17
c92 205 27 1.1226e-16
c93 203 27 8.24397e-17
c94 201 27 1.1226e-16
c95 199 27 1.47899e-17
c96 195 27 1.47899e-17
c97 155 27 1.42959e-16
c98 10 27 1.40799e-17
c99 11 27 1.44349e-16
c100 153 27 1.42959e-16
c101 216 27 1.40799e-17
c102 64 27 1.44349e-16
c103 212 27 9.97196e-17
c104 210 27 9.97196e-17
c105 197 27 1.58499e-17
c106 326 27 3.23999e-18
c107 193 27 1.58499e-17
c108 325 27 3.23999e-18
c109 109 27 6.30198e-17
c110 107 27 6.30198e-17
c111 206 27 6.12598e-17
c112 204 27 8.02596e-17
c113 202 27 6.12598e-17
c114 200 27 8.02596e-17
c115 323 27 3.70198e-17
c116 321 27 3.70198e-17
c117 198 27 7.55907e-17
c118 194 27 7.55907e-17
c119 191 27 2.10199e-17
c120 189 27 2.10199e-17
c121 173 27 1.26499e-17
c122 184 27 1.05821e-16
c123 171 27 1.26499e-17
c124 180 27 1.05821e-16
c125 324 27 4.94098e-17
c126 322 27 4.94098e-17
c127 320 27 2.67999e-18
c128 169 27 1.51099e-17
c129 319 27 2.67999e-18
c130 175 27 1.51099e-17
c131 167 27 1.37899e-17
c132 163 27 1.37899e-17
c133 172 27 8.22296e-17
c134 170 27 8.22296e-17
c135 159 27 1.63299e-17
c136 318 27 3.19999e-18
c137 157 27 1.63299e-17
c138 317 27 3.19999e-18
c139 166 27 7.62606e-17
c140 164 27 6.12607e-17
c141 162 27 7.62606e-17
c142 160 27 6.12607e-17
c143 356 27 3.94304e-17
c144 355 27 2.03004e-17
c145 354 27 3.94304e-17
c146 353 27 2.03004e-17
c147 154 27 8.39596e-17
c148 12 27 1.14349e-16
c149 152 27 8.39596e-17
c150 151 27 1.14349e-16
c151 148 27 1.33799e-17
c152 146 27 1.33799e-17
c153 316 27 2.37999e-18
c154 144 27 1.51099e-17
c155 315 27 2.37999e-18
c156 150 27 1.51099e-17
c157 352 27 2.32404e-17
c158 350 27 3.80801e-17
c159 165 27 1.37899e-17
c160 351 27 2.32404e-17
c161 349 27 3.80801e-17
c162 161 27 1.37899e-17
c163 147 27 8.07997e-17
c164 145 27 8.07997e-17
c165 308 27 3.74099e-17
c166 142 27 1.53299e-17
c167 314 27 3.19999e-18
c168 307 27 3.74099e-17
c169 140 27 1.53299e-17
c170 313 27 3.19999e-18
c171 138 27 1.295e-17
c172 137 27 1.295e-17
c173 124 27 5.89797e-17
c174 122 27 5.89797e-17
c175 312 27 2.67999e-18
c176 134 27 1.51099e-17
c177 311 27 2.67999e-18
c178 136 27 1.51099e-17
c179 185 27 1.37899e-17
c180 181 27 1.37899e-17
c181 128 27 1.63299e-17
c182 310 27 3.19999e-18
c183 126 27 1.63299e-17
c184 309 27 3.19999e-18
c185 114 27 2.30199e-17
c186 306 27 2.40199e-17
c187 112 27 2.30199e-17
c188 304 27 2.40199e-17
c189 119 27 1.11799e-17
c190 117 27 1.11799e-17
c191 305 27 1.51599e-17
c192 303 27 1.51599e-17
c193 115 27 5.29098e-17
c194 116 27 5.29098e-17
c195 13 27 2.03099e-17
c196 14 27 2.03099e-17
c197 110 27 5.11798e-17
c198 15 27 5.11798e-17
c199 16 27 2.59799e-17
c200 103 27 3.99799e-17
c201 108 27 1.39259e-16
c202 106 27 1.39259e-16
c203 105 27 3.44299e-17
c204 17 27 4.68198e-17
c205 104 27 3.44299e-17
c206 102 27 4.68198e-17
c207 18 27 2.74601e-17
c208 302 27 2.74601e-17
c209 95 27 1.37499e-17
c210 93 27 1.37499e-17
c211 101 27 2.11799e-17
c212 100 27 1.74799e-17
c213 99 27 2.11799e-17
c214 98 27 1.74799e-17
c215 301 27 2.57999e-18
c216 91 27 1.62599e-17
c217 300 27 2.57999e-18
c218 97 27 1.62599e-17
c219 89 27 8.24397e-17
c220 87 27 1.1226e-16
c221 85 27 8.24397e-17
c222 83 27 1.1226e-16
c223 20 27 1.47899e-17
c224 80 27 1.47899e-17
c225 94 27 9.97196e-17
c226 92 27 9.97196e-17
c227 21 27 1.58499e-17
c228 299 27 3.23999e-18
c229 78 27 1.58499e-17
c230 298 27 3.23999e-18
c231 88 27 6.12598e-17
c232 86 27 8.02596e-17
c233 84 27 6.12598e-17
c234 82 27 8.02596e-17
c235 296 27 3.70198e-17
c236 294 27 3.70198e-17
c237 22 27 7.55907e-17
c238 79 27 7.55907e-17
c239 76 27 2.10199e-17
c240 74 27 2.10199e-17
c241 60 27 1.26499e-17
c242 70 27 1.05821e-16
c243 58 27 1.26499e-17
c244 66 27 1.05821e-16
c245 297 27 4.94098e-17
c246 295 27 4.94098e-17
c247 293 27 2.67999e-18
c248 56 27 1.51099e-17
c249 292 27 2.67999e-18
c250 62 27 1.51099e-17
c251 54 27 1.37899e-17
c252 52 27 1.37899e-17
c253 59 27 8.22296e-17
c254 57 27 8.22296e-17
c255 48 27 1.63299e-17
c256 291 27 3.19999e-18
c257 46 27 1.63299e-17
c258 290 27 3.19999e-18
c259 23 27 7.62606e-17
c260 24 27 6.12607e-17
c261 51 27 7.62606e-17
c262 49 27 6.12607e-17
c263 348 27 3.94304e-17
c264 347 27 2.03004e-17
c265 346 27 3.94304e-17
c266 345 27 2.03004e-17
c267 42 27 1.33799e-17
c268 40 27 1.33799e-17
c269 289 27 2.37999e-18
c270 38 27 1.51099e-17
c271 288 27 2.37999e-18
c272 44 27 1.51099e-17
c273 344 27 2.32404e-17
c274 342 27 3.80801e-17
c275 53 27 1.37899e-17
c276 343 27 2.32404e-17
c277 341 27 3.80801e-17
c278 50 27 1.37899e-17
c279 41 27 8.07997e-17
c280 39 27 8.07997e-17
c281 336 27 3.74099e-17
c282 36 27 1.53299e-17
c283 287 27 3.19999e-18
c284 335 27 3.74099e-17
c285 34 27 1.53299e-17
c286 286 27 3.19999e-18
c287 32 27 1.295e-17
c288 30 27 1.295e-17
c289 31 27 5.89797e-17
c290 29 27 5.89797e-17
.ends four
.subckt o 1 2 3 4 5
md754 4 7 6 4 penh l=3e-06 w=0.000102 
+ as=4.59e-10 ad=1.258e-09 ps=8.55945e-06 pd=6.84443e-05 
+ nrs=0.0441176 nrd=0.120915 
md755 6 7 4 4 penh l=3e-06 w=0.000102 
+ as=1.258e-09 ad=4.59e-10 ps=6.84443e-05 pd=8.55945e-06 
+ nrs=0.120915 nrd=0.0441176 
md756 4 7 6 4 penh l=3e-06 w=0.0001125 
+ as=5.0625e-10 ad=1.3875e-09 ps=9.44055e-06 pd=7.54901e-05 
+ nrs=0.04 nrd=0.10963 
md757 6 7 4 4 penh l=3e-06 w=0.0001125 
+ as=1.3875e-09 ad=5.0625e-10 ps=7.54901e-05 pd=9.44055e-06 
+ nrs=0.10963 nrd=0.04 
md758 4 6 1 4 penh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.627e-09 ps=2.7e-05 pd=0.000142928 
+ nrs=0.0633802 nrd=0.0579029 
md759 1 6 4 4 penh l=3e-06 w=0.000213 
+ as=2.627e-09 ad=2.8755e-09 ps=0.000142928 pd=2.7e-05 
+ nrs=0.0579029 nrd=0.0633802 
md760 4 6 1 4 penh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.627e-09 ps=2.7e-05 pd=0.000142928 
+ nrs=0.0633802 nrd=0.0579029 
md761 1 6 4 4 penh l=3e-06 w=0.000213 
+ as=2.627e-09 ad=2.8755e-09 ps=0.000142928 pd=2.7e-05 
+ nrs=0.0579029 nrd=0.0633802 
md762 4 6 1 4 penh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.627e-09 ps=2.7e-05 pd=0.000142928 
+ nrs=0.0633802 nrd=0.0579029 
md763 1 6 4 4 penh l=3e-06 w=0.000213 
+ as=2.627e-09 ad=2.8755e-09 ps=0.000142928 pd=2.7e-05 
+ nrs=0.0579029 nrd=0.0633802 
md764 4 6 1 4 penh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.627e-09 ps=2.7e-05 pd=0.000142928 
+ nrs=0.0633802 nrd=0.0579029 
md765 1 6 4 4 penh l=3e-06 w=0.000213 
+ as=2.627e-09 ad=2.8755e-09 ps=0.000142928 pd=2.7e-05 
+ nrs=0.0579029 nrd=0.0633802 
md766 4 5 8 4 penh l=3e-06 w=5.1e-05 
+ as=3.825e-10 ad=6.28999e-10 ps=6.6e-05 pd=3.42222e-05 
+ nrs=0.147059 nrd=0.24183 
md767 7 8 4 4 penh l=3e-06 w=0.000105 
+ as=1.295e-09 ad=7.875e-10 ps=7.04574e-05 pd=0.00012 
+ nrs=0.11746 nrd=0.0714285 
md768 9 5 4 4 penh l=3e-06 w=5.1e-05 
+ as=6.28999e-10 ad=4.545e-10 ps=3.42222e-05 pd=6.9e-05 
+ nrs=0.24183 nrd=0.17474 
md769 10 9 4 4 penh l=3e-06 w=0.0001005 
+ as=1.2395e-09 ad=7.5375e-10 ps=6.74377e-05 pd=0.0001155 
+ nrs=0.12272 nrd=0.0746268 
md770 11 10 4 4 penh l=3e-06 w=0.000102 
+ as=1.258e-09 ad=7.65e-10 ps=6.84443e-05 pd=0.000116641 
+ nrs=0.120915 nrd=0.0735294 
md771 4 10 11 4 penh l=3e-06 w=0.000102 
+ as=7.65e-10 ad=1.258e-09 ps=0.000116641 pd=6.84443e-05 
+ nrs=0.0735294 nrd=0.120915 
md772 4 10 11 4 penh l=3e-06 w=0.0001095 
+ as=8.2125e-10 ad=1.3505e-09 ps=0.000125218 pd=7.34771e-05 
+ nrs=0.0684931 nrd=0.112633 
md773 3 7 6 3 nenh l=3e-06 w=0.00012 
+ as=5.4e-10 ad=1.30558e-09 ps=1.01408e-05 pd=6.68217e-05 
+ nrs=0.0375 nrd=0.0906652 
md774 6 7 3 3 nenh l=3e-06 w=0.00012 
+ as=1.30558e-09 ad=5.4e-10 ps=6.68217e-05 pd=1.01408e-05 
+ nrs=0.0906652 nrd=0.0375 
md775 3 7 6 3 nenh l=3e-06 w=9.3e-05 
+ as=4.185e-10 ad=1.01183e-09 ps=7.85916e-06 pd=5.17868e-05 
+ nrs=0.0483871 nrd=0.116987 
md776 6 7 3 3 nenh l=3e-06 w=9.3e-05 
+ as=1.01183e-09 ad=4.185e-10 ps=5.17868e-05 pd=7.85916e-06 
+ nrs=0.116987 nrd=0.0483871 
md777 3 11 1 3 nenh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.3174e-09 ps=2.7e-05 pd=0.000118608 
+ nrs=0.0633802 nrd=0.051079 
md778 1 11 3 3 nenh l=3e-06 w=0.000213 
+ as=2.3174e-09 ad=2.8755e-09 ps=0.000118608 pd=2.7e-05 
+ nrs=0.051079 nrd=0.0633802 
md779 3 11 1 3 nenh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.3174e-09 ps=2.7e-05 pd=0.000118608 
+ nrs=0.0633802 nrd=0.051079 
md780 1 11 3 3 nenh l=3e-06 w=0.000213 
+ as=2.3174e-09 ad=2.8755e-09 ps=0.000118608 pd=2.7e-05 
+ nrs=0.051079 nrd=0.0633802 
md781 3 11 1 3 nenh l=3e-06 w=0.000213 
+ as=2.8755e-09 ad=2.3174e-09 ps=2.7e-05 pd=0.000118608 
+ nrs=0.0633802 nrd=0.051079 
md782 1 11 3 3 nenh l=3e-06 w=0.000213 
+ as=2.3174e-09 ad=2.8755e-09 ps=0.000118608 pd=2.7e-05 
+ nrs=0.051079 nrd=0.0633802 
md783 3 5 8 3 nenh l=3e-06 w=5.1e-05 
+ as=5.0175e-10 ad=5.54871e-10 ps=7.2e-05 pd=2.83992e-05 
+ nrs=0.192906 nrd=0.21333 
md784 7 8 3 3 nenh l=3e-06 w=0.000105 
+ as=1.14238e-09 ad=7.875e-10 ps=5.84689e-05 pd=0.00012 
+ nrs=0.103618 nrd=0.0714285 
md785 9 5 3 3 nenh l=3e-06 w=5.1e-05 
+ as=5.54871e-10 ad=3.825e-10 ps=2.83992e-05 pd=6.6e-05 
+ nrs=0.21333 nrd=0.147059 
md786 3 9 10 3 nenh l=3e-06 w=0.0001065 
+ as=7.9875e-10 ad=1.1587e-09 ps=0.0001215 pd=5.93042e-05 
+ nrs=0.0704225 nrd=0.102158 
md787 3 10 11 3 nenh l=3e-06 w=9.75e-05 
+ as=5.43934e-10 ad=1.06078e-09 ps=4.56281e-05 pd=5.42926e-05 
+ nrs=0.0572186 nrd=0.111588 
md788 11 10 3 3 nenh l=3e-06 w=0.0001005 
+ as=1.09342e-09 ad=5.6067e-10 ps=5.59631e-05 pd=4.7032e-05 
+ nrs=0.108257 nrd=0.0555106 
md789 11 10 3 3 nenh l=3e-06 w=0.0001065 
+ as=1.1587e-09 ad=5.94144e-10 ps=5.93042e-05 pd=4.98398e-05 
+ nrs=0.102158 nrd=0.0523832 
c291 11 3 1.44725e-16
c292 10 3 4.60348e-17
c293 9 3 5.28303e-17
c294 7 3 8.22997e-17
c295 8 3 5.37903e-17
c296 1 3 1.49951e-15
c297 6 3 1.96039e-16
.ends o
.subckt mcnc#pad 1 2 3 4
c298 1 4 1.049e-18
.ends mcnc#pad
xi#5 1 0 1 3 4 i
xi#4 1 0 1 8 9 i
xi#3 1 0 1 13 14 i
xi#2 1 0 1 18 19 i
xi#1 1 0 1 23 24 i
xi#0 1 0 1 28 29 i
xfour#0 8 3 33 34 35
+ 36 37 38 28 39 40
+ 41 42 43 44 45 46
+ 47 23 48 49 50 51
+ 52 13 18 0 1 four
xo#0 381 1 0 1 42 o
xo#1 388 1 0 1 43 o
xo#2 395 1 0 1 38 o
xo#3 402 1 0 1 45 o
xmcnc#pad#4 0 1 1 1 mcnc#pad
xmcnc#pad#5 0 1 1 0 mcnc#pad
Vshift 4 0 pwl (0 0 8.25e-06 0 8.252e-06 5 8.825e-05 5 
+ 8.8252e-05 0 )
Vexecute 9 0 pwl (0 0 5e-07 0 5.02e-07 5 1e-06 5 
+ 1.002e-06 0 1.5e-06 0 1.502e-06 5 2e-06 5 
+ 2.002e-06 0 2.5e-06 0 2.502e-06 5 3e-06 5 
+ 3.002e-06 0 3.5e-06 0 3.502e-06 5 4e-06 5 
+ 4.002e-06 0 4.5e-06 0 4.502e-06 5 5e-06 5 
+ 5.002e-06 0 5.5e-06 0 5.502e-06 5 6e-06 5 
+ 6.002e-06 0 6.5e-06 0 6.502e-06 5 7e-06 5 
+ 7.002e-06 0 7.5e-06 0 7.502e-06 5 8e-06 5 
+ 8.002e-06 0 8.5e-06 0 8.502e-06 5 9e-06 5 
+ 9.002e-06 0 9.5e-06 0 9.502e-06 5 1e-05 5 
+ 1.0002e-05 0 1.05e-05 0 1.0502e-05 5 1.1e-05 5 
+ 1.1002e-05 0 1.15e-05 0 1.1502e-05 5 1.2e-05 5 
+ 1.2002e-05 0 1.25e-05 0 1.2502e-05 5 1.3e-05 5 
+ 1.3002e-05 0 1.35e-05 0 1.3502e-05 5 1.4e-05 5 
+ 1.4002e-05 0 1.45e-05 0 1.4502e-05 5 1.5e-05 5 
+ 1.5002e-05 0 1.55e-05 0 1.5502e-05 5 1.6e-05 5 
+ 1.6002e-05 0 1.65e-05 0 1.6502e-05 5 1.7e-05 5 
+ 1.7002e-05 0 1.75e-05 0 1.7502e-05 5 1.8e-05 5 
+ 1.8002e-05 0 1.85e-05 0 1.8502e-05 5 1.9e-05 5 
+ 1.9002e-05 0 1.95e-05 0 1.9502e-05 5 2e-05 5 
+ 2.0002e-05 0 2.05e-05 0 2.0502e-05 5 2.1e-05 5 
+ 2.1002e-05 0 2.15e-05 0 2.1502e-05 5 2.2e-05 5 
+ 2.2002e-05 0 2.25e-05 0 2.2502e-05 5 2.3e-05 5 
+ 2.3002e-05 0 2.35e-05 0 2.3502e-05 5 2.4e-05 5 
+ 2.4002e-05 0 )
Vx1in 24 0 pwl (0 0 1.25e-06 0 1.252e-06 5 2.25e-06 5 
+ 2.252e-06 0 3.25e-06 0 3.252e-06 5 4.25e-06 5 
+ 4.252e-06 0 5.25e-06 0 5.252e-06 5 6.25e-06 5 
+ 6.252e-06 0 7.25e-06 0 7.252e-06 5 8.25e-06 5 
+ 8.252e-06 0 1.425e-05 0 1.4252e-05 5 2.025e-05 5 
+ 2.0252e-05 0 2.125e-05 0 2.1252e-05 5 2.225e-05 5 
+ 2.2252e-05 0 2.325e-05 0 2.3252e-05 5 2.425e-05 5 
+ 2.4252e-05 0 )
Vx2in 29 0 pwl (0 0 1.25e-06 0 1.252e-06 5 2.25e-06 5 
+ 2.252e-06 0 3.25e-06 0 3.252e-06 5 4.25e-06 5 
+ 4.252e-06 0 5.25e-06 0 5.252e-06 5 6.25e-06 5 
+ 6.252e-06 0 7.25e-06 0 7.252e-06 5 8.25e-06 5 
+ 8.252e-06 0 1.325e-05 0 1.3252e-05 5 1.425e-05 5 
+ 1.4252e-05 0 1.525e-05 0 1.5252e-05 5 2.025e-05 5 
+ 2.0252e-05 0 2.225e-05 0 2.2252e-05 5 2.425e-05 5 
+ 2.4252e-05 0 )
Vy1in 19 0 pwl (0 0 1.25e-06 0 1.252e-06 5 2.25e-06 5 
+ 2.252e-06 0 3.25e-06 0 3.252e-06 5 4.25e-06 5 
+ 4.252e-06 0 5.25e-06 0 5.252e-06 5 6.25e-06 5 
+ 6.252e-06 0 7.25e-06 0 7.252e-06 5 8.25e-06 5 
+ 8.252e-06 0 1.025e-05 0 1.0252e-05 5 1.225e-05 5 
+ 1.2252e-05 0 1.625e-05 0 1.6252e-05 5 2.025e-05 5 
+ 2.0252e-05 0 2.125e-05 0 2.1252e-05 5 2.225e-05 5 
+ 2.2252e-05 0 2.325e-05 0 2.3252e-05 5 2.425e-05 5 
+ 2.4252e-05 0 )
Vy2in 14 0 pwl (0 0 1.25e-06 0 1.252e-06 5 2.25e-06 5 
+ 2.252e-06 0 3.25e-06 0 3.252e-06 5 4.25e-06 5 
+ 4.252e-06 0 5.25e-06 0 5.252e-06 5 6.25e-06 5 
+ 6.252e-06 0 7.25e-06 0 7.252e-06 5 8.25e-06 5 
+ 8.252e-06 0 9.25e-06 0 9.252e-06 5 1.025e-05 5 
+ 1.0252e-05 0 1.125e-05 0 1.1252e-05 5 1.225e-05 5 
+ 1.2252e-05 0 1.625e-05 0 1.6252e-05 5 2.025e-05 5 
+ 2.0252e-05 0 2.225e-05 0 2.2252e-05 5 2.425e-05 5 
+ 2.4252e-05 0 )
VVDD 1 0 5
.temp 75 
*.print TRAN v(9) v(4) v(23) v(46) v(35) v(37) 
+v(49) v(48) v(50) v(40) v(41) v(3) 
+v(34) v(33) v(36) v(39) v(24) v(29) 
+v(19) v(14) v(402) v(388) 
.options limpts=50000 itl5=50000
*.TRAN 1e-07 2.4e-05
.op
.end
