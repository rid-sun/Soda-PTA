HYBRID VOLTAGE REFERENCE 2000.12.18 Y.I
*.OP
*.TRAN 1 50 0 1
VCC 50 0 DC 5.0
R1 6 1 948.0
R2 6 2 2.844K
R3 3 0 362.0
R5 50 7 3.100K
R6 50 4 3.28K
R7 5 6 3.2K
R8 1 8 362.0
Q1 1 1 0 QNPN
Q2 2 8 3 QNPN 3.33
Q3 4 2 0 QNPN
Q4 50 4 6 QNPN 3.33
Q5 4 7 5 QNPN
Q6 5 5 0 QNPN
Q7 7 8 0 QNPN
Q8 9 5 0 QNPN
Q9 7 7 9 QNPN
*Q10 7 7 6 QNPN
.MODEL QNPN NPN (IS=1.0E-16 BF=100 BR=1 VAF=0)
*.PRINT TRAN V(100) V(101) I(VCC)
*.PRINT TRAN V(1) V(2) V(3) V(4) V(5) V(6) V(7) V(8) V(9) V(50)
*.END

.OPTIONS DELMAX=1000ns
.op
*.pstran convval=1.0e-05 initstep=1.0e-05 minstep=1.0e-09 maxstep=1.0e+6 tau=1.0e-05 vbe0=0.0 kvgs0=0.0  tauramp=0.0
.end 