TADEGLOW6TR CKT
VCC 1 0 DC 12.0
RT1C 1 2 2.7K
RT1B 4 5 5.0K
RT2CD 3 5 15.0K
RT2C 1 5 2.7K
RT3CD 8 6 15.0K
RT3C 1 8 1.0K
RT3B 9 10 15.0K
RT34E 11 0 50.0
RT4C 1 10 3.0K
RT4B1 1 12 11.0K
RT4B2 12 0 1.0K
RT5C 1 13 11.0K
RT5CD 13 7 15.0K
RT5B 14 15 15.0K
RT56E 16 0 50.0
RT6C 1 15 3.0K
RT6B1 1 17 11.0K
RT6B2 17 0 1.0K
DT1 2 3 DIODE
DT3 6 5 DIODE
DT5 7 5 DIODE
QT1 2 4 0 QNPN
QT2 5 5 0 QNPN
QT3 8 9 11 QNPN
QT4 10 12 11 QNPN
QT5 13 14 16 QNPN
QT6 15 17 16 QNPN
.MODEL DIODE D (IS=1.0E-14)
.MODEL QNPN NPN (IS=1.0E-14 BF=100 VA=50)
*.END

.OPTIONS DELMAX=1000ns
.op
*.gmin
.end 